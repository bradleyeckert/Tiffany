library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

-- Single-port synchronous-read ROM

ENTITY ROM32 IS
generic (
  Size:  integer := 10                          -- log2 (cells)
);
port (
  clk:    in  std_logic;                        -- System clock
  addr:   in  std_logic_vector(Size-1 downto 0);
  data_o: out std_logic_vector(31 downto 0)     -- read data
);
END ROM32;

ARCHITECTURE RTL OF ROM32 IS
signal address: integer range 0 to 2**Size-1;
begin
address <= to_integer(unsigned(addr));

process (clk) begin
  if rising_edge(clk) then
    case address is
      when   0 => data_o <= x"54000281";
      when   1 => data_o <= x"54000284";
      when   2 => data_o <= x"54000000";
      when   3 => data_o <= x"D090C220";
      when   4 => data_o <= x"9FB08800";
      when   5 => data_o <= x"3FB08800";
      when   6 => data_o <= x"5FB08800";
      when   7 => data_o <= x"05FB8328";
      when   8 => data_o <= x"9FB08800";
      when   9 => data_o <= x"05FD8328";
      when  10 => data_o <= x"3FB08800";
      when  11 => data_o <= x"D0908800";
      when  12 => data_o <= x"D09D0220";
      when  13 => data_o <= x"D21D0220";
      when  14 => data_o <= x"10408800";
      when  15 => data_o <= x"7FC2BC08";
      when  16 => data_o <= x"F1FF0A08";
      when  17 => data_o <= x"F3908800";
      when  18 => data_o <= x"F3B08800";
      when  19 => data_o <= x"F0AF1FF0";
      when  20 => data_o <= x"7DF08800";
      when  21 => data_o <= x"28AF0AF0";
      when  22 => data_o <= x"7FC08800";
      when  23 => data_o <= x"28A4BC7C";
      when  24 => data_o <= x"F12F1F08";
      when  25 => data_o <= x"EFB08800";
      when  26 => data_o <= x"E7908800";
      when  27 => data_o <= x"7FC2BC7C";
      when  28 => data_o <= x"7FC2BC2A";
      when  29 => data_o <= x"7DFE7928";
      when  30 => data_o <= x"2950001B";
      when  31 => data_o <= x"EFBEC220";
      when  32 => data_o <= x"07A08800";
      when  33 => data_o <= x"04220000";
      when  34 => data_o <= x"07005BD2";
      when  35 => data_o <= x"05B08800";
      when  36 => data_o <= x"90220000";
      when  37 => data_o <= x"6E408800";
      when  38 => data_o <= x"6E490220";
      when  39 => data_o <= x"92408800";
      when  40 => data_o <= x"D09B0220";
      when  41 => data_o <= x"24927D03";
      when  42 => data_o <= x"D1308800";
      when  43 => data_o <= x"9BCBBC08";
      when  44 => data_o <= x"9E7EC220";
      when  45 => data_o <= x"C3424800";
      when  46 => data_o <= x"08800000";
      when  47 => data_o <= x"D3CD13D2";
      when  48 => data_o <= x"7C220000";
      when  49 => data_o <= x"7DFF0A0C";
      when  50 => data_o <= x"F0A8C220";
      when  51 => data_o <= x"D1FD0928";
      when  52 => data_o <= x"E64C3B26";
      when  53 => data_o <= x"EC220000";
      when  54 => data_o <= x"C1500033";
      when  55 => data_o <= x"08800000";
      when  56 => data_o <= x"38220000";
      when  57 => data_o <= x"F4000004";
      when  58 => data_o <= x"66E08800";
      when  59 => data_o <= x"F4000008";
      when  60 => data_o <= x"66E08800";
      when  61 => data_o <= x"F400000C";
      when  62 => data_o <= x"A6EF4008";
      when  63 => data_o <= x"67424350";
      when  64 => data_o <= x"50220000";
      when  65 => data_o <= x"044119B8";
      when  66 => data_o <= x"F3B08800";
      when  67 => data_o <= x"F400000A";
      when  68 => data_o <= x"F4000DE7";
      when  69 => data_o <= x"D27EC220";
      when  70 => data_o <= x"F4000010";
      when  71 => data_o <= x"F4000DE7";
      when  72 => data_o <= x"D27EC220";
      when  73 => data_o <= x"B8800000";
      when  74 => data_o <= x"F4FFFFFF";
      when  75 => data_o <= x"4C220000";
      when  76 => data_o <= x"E79D0320";
      when  77 => data_o <= x"C3BEFB08";
      when  78 => data_o <= x"EFCD0928";
      when  79 => data_o <= x"87C7FC7C";
      when  80 => data_o <= x"7C220000";
      when  81 => data_o <= x"28A24AE4";
      when  82 => data_o <= x"E4320000";
      when  83 => data_o <= x"C3B7DF7E";
      when  84 => data_o <= x"EFBEE17E";
      when  85 => data_o <= x"2BC2B90C";
      when  86 => data_o <= x"4B90FC7C";
      when  87 => data_o <= x"F2C6C800";
      when  88 => data_o <= x"C3B7C220";
      when  89 => data_o <= x"ECAECAEC";
      when  90 => data_o <= x"85F08800";
      when  91 => data_o <= x"F400000C";
      when  92 => data_o <= x"46E08800";
      when  93 => data_o <= x"28AECAEC";
      when  94 => data_o <= x"7C220000";
      when  95 => data_o <= x"E796E420";
      when  96 => data_o <= x"EBB08800";
      when  97 => data_o <= x"EFB2A17E";
      when  98 => data_o <= x"28AD09D0";
      when  99 => data_o <= x"C3B7C220";
      when 100 => data_o <= x"7E17C220";
      when 101 => data_o <= x"281383F7";
      when 102 => data_o <= x"05F0CAD0";
      when 103 => data_o <= x"4DF08800";
      when 104 => data_o <= x"D090CCF5";
      when 105 => data_o <= x"4F427408";
      when 106 => data_o <= x"F1500068";
      when 107 => data_o <= x"E796EC20";
      when 108 => data_o <= x"EB4243B2";
      when 109 => data_o <= x"EEC08800";
      when 110 => data_o <= x"F150006B";
      when 111 => data_o <= x"D09D0800";
      when 112 => data_o <= x"C1500074";
      when 113 => data_o <= x"D09F1FF0";
      when 114 => data_o <= x"98A9DFA0";
      when 115 => data_o <= x"2BBEFB08";
      when 116 => data_o <= x"EFBEC220";
      when 117 => data_o <= x"D09D0800";
      when 118 => data_o <= x"C150007A";
      when 119 => data_o <= x"D09F1FF0";
      when 120 => data_o <= x"38A3DFA0";
      when 121 => data_o <= x"2BBEFB08";
      when 122 => data_o <= x"EFBEC220";
      when 123 => data_o <= x"D09D0800";
      when 124 => data_o <= x"C1500084";
      when 125 => data_o <= x"2417C3F0";
      when 126 => data_o <= x"483F0AD0";
      when 127 => data_o <= x"24800000";
      when 128 => data_o <= x"7F4274F0";
      when 129 => data_o <= x"D09D3CE4";
      when 130 => data_o <= x"DB93FB28";
      when 131 => data_o <= x"27054080";
      when 132 => data_o <= x"EFBEC220";
      when 133 => data_o <= x"7F9E5D68";
      when 134 => data_o <= x"E9500089";
      when 135 => data_o <= x"29D0007B";
      when 136 => data_o <= x"5400008A";
      when 137 => data_o <= x"29D00075";
      when 138 => data_o <= x"08800000";
      when 139 => data_o <= x"E7A54090";
      when 140 => data_o <= x"F34249F0";
      when 141 => data_o <= x"7FC20000";
      when 142 => data_o <= x"4BC3E828";
      when 143 => data_o <= x"EFBEC220";
      when 144 => data_o <= x"EFBEC220";
      when 145 => data_o <= x"07AEFB08";
      when 146 => data_o <= x"E797402F";
      when 147 => data_o <= x"F4000003";
      when 148 => data_o <= x"4FA54097";
      when 149 => data_o <= x"F4000000";
      when 150 => data_o <= x"5400008B";
      when 151 => data_o <= x"0416DF50";
      when 152 => data_o <= x"534249F0";
      when 153 => data_o <= x"4BC9E828";
      when 154 => data_o <= x"EFBEC220";
      when 155 => data_o <= x"D09D30EE";
      when 156 => data_o <= x"F400003F";
      when 157 => data_o <= x"4F427C20";
      when 158 => data_o <= x"128F3B08";
      when 159 => data_o <= x"08800000";
      when 160 => data_o <= x"D09D30EE";
      when 161 => data_o <= x"F400003F";
      when 162 => data_o <= x"4F427C20";
      when 163 => data_o <= x"728F3B08";
      when 164 => data_o <= x"08800000";
      when 165 => data_o <= x"0416FD1F";
      when 166 => data_o <= x"D0800000";
      when 167 => data_o <= x"7C47CC20";
      when 168 => data_o <= x"E392837C";
      when 169 => data_o <= x"E0920000";
      when 170 => data_o <= x"28A24800";
      when 171 => data_o <= x"C15000A7";
      when 172 => data_o <= x"EDF7FB28";
      when 173 => data_o <= x"2BC08800";
      when 174 => data_o <= x"E79D090C";
      when 175 => data_o <= x"EF8540BE";
      when 176 => data_o <= x"F400001F";
      when 177 => data_o <= x"D1C10800";
      when 178 => data_o <= x"7DFF0CF0";
      when 179 => data_o <= x"338540B9";
      when 180 => data_o <= x"052D090C";
      when 181 => data_o <= x"EC800000";
      when 182 => data_o <= x"E12D090C";
      when 183 => data_o <= x"04CD14EC";
      when 184 => data_o <= x"540000BB";
      when 185 => data_o <= x"4B4243F4";
      when 186 => data_o <= x"13B20000";
      when 187 => data_o <= x"28A24800";
      when 188 => data_o <= x"C15000B2";
      when 189 => data_o <= x"EFBF0CD2";
      when 190 => data_o <= x"EFBEFD00";
      when 191 => data_o <= x"D0108800";
      when 192 => data_o <= x"E796DFE4";
      when 193 => data_o <= x"7DD0002D";
      when 194 => data_o <= x"7DD00036";
      when 195 => data_o <= x"29D000AE";
      when 196 => data_o <= x"F0AB0800";
      when 197 => data_o <= x"E95000C7";
      when 198 => data_o <= x"D0920000";
      when 199 => data_o <= x"F0AB0800";
      when 200 => data_o <= x"E95000CA";
      when 201 => data_o <= x"D0920000";
      when 202 => data_o <= x"08800000";
      when 203 => data_o <= x"05FE796C";
      when 204 => data_o <= x"7C17DD2D";
      when 205 => data_o <= x"7DD00036";
      when 206 => data_o <= x"29D000AE";
      when 207 => data_o <= x"F0AB0800";
      when 208 => data_o <= x"E95000D2";
      when 209 => data_o <= x"D0920000";
      when 210 => data_o <= x"F0AB0800";
      when 211 => data_o <= x"E95000D9";
      when 212 => data_o <= x"D09E4800";
      when 213 => data_o <= x"E95000D9";
      when 214 => data_o <= x"49FF0AF0";
      when 215 => data_o <= x"D090FCD0";
      when 216 => data_o <= x"27420000";
      when 217 => data_o <= x"2BB08800";
      when 218 => data_o <= x"06C05F20";
      when 219 => data_o <= x"E95000DE";
      when 220 => data_o <= x"D097DD33";
      when 221 => data_o <= x"28800000";
      when 222 => data_o <= x"7C1B0800";
      when 223 => data_o <= x"E95000E1";
      when 224 => data_o <= x"48320000";
      when 225 => data_o <= x"29D000AE";
      when 226 => data_o <= x"2BA540E4";
      when 227 => data_o <= x"F3427C20";
      when 228 => data_o <= x"08800000";
      when 229 => data_o <= x"E6CF15DA";
      when 230 => data_o <= x"740000E5";
      when 231 => data_o <= x"EC220000";
      when 232 => data_o <= x"740000E5";
      when 233 => data_o <= x"F3B08800";
      when 234 => data_o <= x"E797406B";
      when 235 => data_o <= x"EBC20000";
      when 236 => data_o <= x"EC220000";
      when 237 => data_o <= x"E79F1D6B";
      when 238 => data_o <= x"EBC20000";
      when 239 => data_o <= x"EC220000";
      when 240 => data_o <= x"E7974068";
      when 241 => data_o <= x"EBC20000";
      when 242 => data_o <= x"EC220000";
      when 243 => data_o <= x"E79F1D68";
      when 244 => data_o <= x"EBC20000";
      when 245 => data_o <= x"EC220000";
      when 246 => data_o <= x"7FC483F0";
      when 247 => data_o <= x"2B424308";
      when 248 => data_o <= x"E742437C";
      when 249 => data_o <= x"D090CA20";
      when 250 => data_o <= x"54000068";
      when 251 => data_o <= x"740000A5";
      when 252 => data_o <= x"EC220000";
      when 253 => data_o <= x"E796EC7C";
      when 254 => data_o <= x"7400002D";
      when 255 => data_o <= x"F1D0002D";
      when 256 => data_o <= x"740000A5";
      when 257 => data_o <= x"2BA54103";
      when 258 => data_o <= x"74000033";
      when 259 => data_o <= x"08800000";
      when 260 => data_o <= x"7DD000FD";
      when 261 => data_o <= x"295000DA";
      when 262 => data_o <= x"74000104";
      when 263 => data_o <= x"F3B08800";
      when 264 => data_o <= x"34000001";
      when 265 => data_o <= x"54000109";
      when 266 => data_o <= x"08800000";
      when 267 => data_o <= x"F3D00000";
      when 268 => data_o <= x"D1F20000";
      when 269 => data_o <= x"E7A54117";
      when 270 => data_o <= x"F34274F0";
      when 271 => data_o <= x"38A6FD07";
      when 272 => data_o <= x"D0800000";
      when 273 => data_o <= x"25F07D01";
      when 274 => data_o <= x"4F427DED";
      when 275 => data_o <= x"94B88320";
      when 276 => data_o <= x"4FC71B28";
      when 277 => data_o <= x"C1500111";
      when 278 => data_o <= x"EDF5410D";
      when 279 => data_o <= x"EFB2B408";
      when 280 => data_o <= x"E5FF4004";
      when 281 => data_o <= x"65FF4DEB";
      when 282 => data_o <= x"D2E7FD00";
      when 283 => data_o <= x"47D00DEB";
      when 284 => data_o <= x"D27EDD30";
      when 285 => data_o <= x"2BD00DEB";
      when 286 => data_o <= x"D27ECAEC";
      when 287 => data_o <= x"2816C220";
      when 288 => data_o <= x"07AEC220";
      when 289 => data_o <= x"F4000DEB";
      when 290 => data_o <= x"D2EBCA20";
      when 291 => data_o <= x"F4000DEB";
      when 292 => data_o <= x"D27ECAF0";
      when 293 => data_o <= x"7F7EFCEC";
      when 294 => data_o <= x"28AF0220";
      when 295 => data_o <= x"08800000";
      when 296 => data_o <= x"04D00002";
      when 297 => data_o <= x"08800000";
      when 298 => data_o <= x"F4000021";
      when 299 => data_o <= x"740000FB";
      when 300 => data_o <= x"74000128";
      when 301 => data_o <= x"0C800000";
      when 302 => data_o <= x"74000127";
      when 303 => data_o <= x"05D00128";
      when 304 => data_o <= x"7400006B";
      when 305 => data_o <= x"E950012E";
      when 306 => data_o <= x"EC220000";
      when 307 => data_o <= x"F3D0FFFF";
      when 308 => data_o <= x"4C334000";
      when 309 => data_o <= x"08800000";
      when 310 => data_o <= x"74000133";
      when 311 => data_o <= x"EC220000";
      when 312 => data_o <= x"74000127";
      when 313 => data_o <= x"F4060000";
      when 314 => data_o <= x"34000000";
      when 315 => data_o <= x"E9500138";
      when 316 => data_o <= x"F4010000";
      when 317 => data_o <= x"54000136";
      when 318 => data_o <= x"54000162";
      when 319 => data_o <= x"3950013E";
      when 320 => data_o <= x"040A0D02";
      when 321 => data_o <= x"4A325B1B";
      when 322 => data_o <= x"F4000500";
      when 323 => data_o <= x"5400013F";
      when 324 => data_o <= x"F4000503";
      when 325 => data_o <= x"5400013F";
      when 326 => data_o <= x"F4000000";
      when 327 => data_o <= x"34000000";
      when 328 => data_o <= x"54000127";
      when 329 => data_o <= x"74000146";
      when 330 => data_o <= x"E9500149";
      when 331 => data_o <= x"F4020000";
      when 332 => data_o <= x"34000000";
      when 333 => data_o <= x"08800000";
      when 334 => data_o <= x"000004E0";
      when 335 => data_o <= x"00000508";
      when 336 => data_o <= x"00000510";
      when 337 => data_o <= x"00000518";
      when 338 => data_o <= x"00000524";
      when 339 => data_o <= x"F4000538";
      when 340 => data_o <= x"F4000DCF";
      when 341 => data_o <= x"D27EC220";
      when 342 => data_o <= x"104F4DCF";
      when 343 => data_o <= x"D2E0EE7E";
      when 344 => data_o <= x"F4000000";
      when 345 => data_o <= x"54000156";
      when 346 => data_o <= x"F4000001";
      when 347 => data_o <= x"54000156";
      when 348 => data_o <= x"F4000002";
      when 349 => data_o <= x"54000156";
      when 350 => data_o <= x"F4000003";
      when 351 => data_o <= x"54000156";
      when 352 => data_o <= x"F4000004";
      when 353 => data_o <= x"54000156";
      when 354 => data_o <= x"07AEFB08";
      when 355 => data_o <= x"D0920000";
      when 356 => data_o <= x"25F38800";
      when 357 => data_o <= x"74000158";
      when 358 => data_o <= x"2B054164";
      when 359 => data_o <= x"EFB08800";
      when 360 => data_o <= x"F4000020";
      when 361 => data_o <= x"54000158";
      when 362 => data_o <= x"C3B08800";
      when 363 => data_o <= x"74000168";
      when 364 => data_o <= x"D09D0800";
      when 365 => data_o <= x"5400016A";
      when 366 => data_o <= x"08800000";
      when 367 => data_o <= x"07D00009";
      when 368 => data_o <= x"D03B3D06";
      when 369 => data_o <= x"D130FD37";
      when 370 => data_o <= x"0C220000";
      when 371 => data_o <= x"F4000CCB";
      when 372 => data_o <= x"D3D00D97";
      when 373 => data_o <= x"D27EC220";
      when 374 => data_o <= x"F4000D97";
      when 375 => data_o <= x"D017EED0";
      when 376 => data_o <= x"27404A9C";
      when 377 => data_o <= x"ECFEC220";
      when 378 => data_o <= x"07D00DE7";
      when 379 => data_o <= x"D2E7C800";
      when 380 => data_o <= x"E9500183";
      when 381 => data_o <= x"F4000000";
      when 382 => data_o <= x"49D000AE";
      when 383 => data_o <= x"2BC7DDAE";
      when 384 => data_o <= x"F1D0016F";
      when 385 => data_o <= x"74000176";
      when 386 => data_o <= x"28220000";
      when 387 => data_o <= x"29D000AE";
      when 388 => data_o <= x"F1D0016F";
      when 389 => data_o <= x"74000176";
      when 390 => data_o <= x"0416C220";
      when 391 => data_o <= x"7400017A";
      when 392 => data_o <= x"E797402F";
      when 393 => data_o <= x"93A54187";
      when 394 => data_o <= x"08800000";
      when 395 => data_o <= x"B3A5418E";
      when 396 => data_o <= x"F400002D";
      when 397 => data_o <= x"74000176";
      when 398 => data_o <= x"08800000";
      when 399 => data_o <= x"EFBF4D97";
      when 400 => data_o <= x"D2EF4CCB";
      when 401 => data_o <= x"D39D090E";
      when 402 => data_o <= x"E7424320";
      when 403 => data_o <= x"7400016A";
      when 404 => data_o <= x"5400013E";
      when 405 => data_o <= x"7C17DD36";
      when 406 => data_o <= x"74000173";
      when 407 => data_o <= x"74000187";
      when 408 => data_o <= x"29D0018B";
      when 409 => data_o <= x"7400018F";
      when 410 => data_o <= x"29500192";
      when 411 => data_o <= x"F4000000";
      when 412 => data_o <= x"F1500195";
      when 413 => data_o <= x"7DD00022";
      when 414 => data_o <= x"29500195";
      when 415 => data_o <= x"F4000000";
      when 416 => data_o <= x"74000195";
      when 417 => data_o <= x"54000168";
      when 418 => data_o <= x"F4000000";
      when 419 => data_o <= x"5400019F";
      when 420 => data_o <= x"F4000DE7";
      when 421 => data_o <= x"D2EF400A";
      when 422 => data_o <= x"6FA541A8";
      when 423 => data_o <= x"540001A2";
      when 424 => data_o <= x"74000022";
      when 425 => data_o <= x"5400019F";
      when 426 => data_o <= x"B95001A4";
      when 427 => data_o <= x"74000173";
      when 428 => data_o <= x"D0920000";
      when 429 => data_o <= x"7DD0017A";
      when 430 => data_o <= x"28920000";
      when 431 => data_o <= x"C15001AD";
      when 432 => data_o <= x"EDD00187";
      when 433 => data_o <= x"5400018F";
      when 434 => data_o <= x"F4000DE7";
      when 435 => data_o <= x"D2E7DD46";
      when 436 => data_o <= x"F4000000";
      when 437 => data_o <= x"F1D001AB";
      when 438 => data_o <= x"2BD00DE7";
      when 439 => data_o <= x"D27EC800";
      when 440 => data_o <= x"7400013E";
      when 441 => data_o <= x"54000168";
      when 442 => data_o <= x"7C104A0C";
      when 443 => data_o <= x"7C800000";
      when 444 => data_o <= x"0526C800";
      when 445 => data_o <= x"E95001DE";
      when 446 => data_o <= x"74000127";
      when 447 => data_o <= x"7400015E";
      when 448 => data_o <= x"E95001BE";
      when 449 => data_o <= x"74000160";
      when 450 => data_o <= x"07D0000D";
      when 451 => data_o <= x"6E420000";
      when 452 => data_o <= x"E95001C7";
      when 453 => data_o <= x"ECAEFCD0";
      when 454 => data_o <= x"24308800";
      when 455 => data_o <= x"07D00008";
      when 456 => data_o <= x"6E420000";
      when 457 => data_o <= x"E95001D3";
      when 458 => data_o <= x"EF9E5B20";
      when 459 => data_o <= x"E95001D2";
      when 460 => data_o <= x"D09D0800";
      when 461 => data_o <= x"540001D0";
      when 462 => data_o <= x"445B1B07";
      when 463 => data_o <= x"445B1B20";
      when 464 => data_o <= x"F4000738";
      when 465 => data_o <= x"39D0013E";
      when 466 => data_o <= x"540001DD";
      when 467 => data_o <= x"07D00020";
      when 468 => data_o <= x"D090C800";
      when 469 => data_o <= x"C15001DC";
      when 470 => data_o <= x"EFD00DB1";
      when 471 => data_o <= x"D3690800";
      when 472 => data_o <= x"E95001DA";
      when 473 => data_o <= x"05D00158";
      when 474 => data_o <= x"F0F20000";
      when 475 => data_o <= x"540001DD";
      when 476 => data_o <= x"EFB20000";
      when 477 => data_o <= x"540001BC";
      when 478 => data_o <= x"2BBF3427";
      when 479 => data_o <= x"08800000";
      when 480 => data_o <= x"9FB08800";
      when 481 => data_o <= x"7F4F40FF";
      when 482 => data_o <= x"4D2F4003";
      when 483 => data_o <= x"4C410420";
      when 484 => data_o <= x"7400009B";
      when 485 => data_o <= x"D0AF4003";
      when 486 => data_o <= x"D139FB08";
      when 487 => data_o <= x"D0920000";
      when 488 => data_o <= x"7F9DB920";
      when 489 => data_o <= x"740001E1";
      when 490 => data_o <= x"27C27C28";
      when 491 => data_o <= x"270541E8";
      when 492 => data_o <= x"EFBEC220";
      when 493 => data_o <= x"F4000000";
      when 494 => data_o <= x"F4000D9C";
      when 495 => data_o <= x"D0FEC220";
      when 496 => data_o <= x"F4000001";
      when 497 => data_o <= x"F4000D9C";
      when 498 => data_o <= x"D0FEC220";
      when 499 => data_o <= x"F4000D9C";
      when 500 => data_o <= x"D3620000";
      when 501 => data_o <= x"E95001F8";
      when 502 => data_o <= x"F4000DDF";
      when 503 => data_o <= x"D0220000";
      when 504 => data_o <= x"F4000DDB";
      when 505 => data_o <= x"D0220000";
      when 506 => data_o <= x"05FB8800";
      when 507 => data_o <= x"740001E0";
      when 508 => data_o <= x"F4000004";
      when 509 => data_o <= x"29500007";
      when 510 => data_o <= x"F4000DDF";
      when 511 => data_o <= x"D15001FA";
      when 512 => data_o <= x"F4000DE3";
      when 513 => data_o <= x"D15001FA";
      when 514 => data_o <= x"F4000DDB";
      when 515 => data_o <= x"D017EE9C";
      when 516 => data_o <= x"EFD00004";
      when 517 => data_o <= x"29500007";
      when 518 => data_o <= x"F4000D9C";
      when 519 => data_o <= x"D3620000";
      when 520 => data_o <= x"E950020A";
      when 521 => data_o <= x"540001FE";
      when 522 => data_o <= x"54000202";
      when 523 => data_o <= x"05FB8800";
      when 524 => data_o <= x"740001E1";
      when 525 => data_o <= x"4AE24A9C";
      when 526 => data_o <= x"EC220000";
      when 527 => data_o <= x"F4000DDF";
      when 528 => data_o <= x"D150020B";
      when 529 => data_o <= x"F4000DE3";
      when 530 => data_o <= x"D150020B";
      when 531 => data_o <= x"F4000DDB";
      when 532 => data_o <= x"D017EE3C";
      when 533 => data_o <= x"EFD00001";
      when 534 => data_o <= x"29500007";
      when 535 => data_o <= x"F4000D9C";
      when 536 => data_o <= x"D3620000";
      when 537 => data_o <= x"E950021B";
      when 538 => data_o <= x"5400020F";
      when 539 => data_o <= x"54000213";
      when 540 => data_o <= x"E7D00DDB";
      when 541 => data_o <= x"D2E6D308";
      when 542 => data_o <= x"F4000DDF";
      when 543 => data_o <= x"D2EF3D00";
      when 544 => data_o <= x"D1D001FE";
      when 545 => data_o <= x"06E90800";
      when 546 => data_o <= x"7400021C";
      when 547 => data_o <= x"E9500225";
      when 548 => data_o <= x"85500221";
      when 549 => data_o <= x"041741FE";
      when 550 => data_o <= x"06E92420";
      when 551 => data_o <= x"7400021C";
      when 552 => data_o <= x"E950022B";
      when 553 => data_o <= x"99D001FE";
      when 554 => data_o <= x"54000226";
      when 555 => data_o <= x"08800000";
      when 556 => data_o <= x"F4000DC7";
      when 557 => data_o <= x"D2EF4DBF";
      when 558 => data_o <= x"D27EC800";
      when 559 => data_o <= x"F4000D97";
      when 560 => data_o <= x"D3D000CC";
      when 561 => data_o <= x"74000091";
      when 562 => data_o <= x"F4000000";
      when 563 => data_o <= x"A4800000";
      when 564 => data_o <= x"7400021E";
      when 565 => data_o <= x"7F42520C";
      when 566 => data_o <= x"514F39F0";
      when 567 => data_o <= x"740001E0";
      when 568 => data_o <= x"2BC90800";
      when 569 => data_o <= x"E9500234";
      when 570 => data_o <= x"EC220000";
      when 571 => data_o <= x"54000240";
      when 572 => data_o <= x"6C65480C";
      when 573 => data_o <= x"57206F6C";
      when 574 => data_o <= x"646C726F";
      when 575 => data_o <= x"FFFFFF21";
      when 576 => data_o <= x"F40008F0";
      when 577 => data_o <= x"39D0013E";
      when 578 => data_o <= x"7400015A";
      when 579 => data_o <= x"F400000A";
      when 580 => data_o <= x"F4000000";
      when 581 => data_o <= x"F3425F7C";
      when 582 => data_o <= x"49D001A4";
      when 583 => data_o <= x"74000051";
      when 584 => data_o <= x"54000246";
      when 585 => data_o <= x"5400015A";
      when 586 => data_o <= x"00000003";
      when 587 => data_o <= x"FFFFF204";
      when 588 => data_o <= x"FFFFF200";
      when 589 => data_o <= x"FFFFF1F0";
      when 590 => data_o <= x"FFFFF100";
      when 591 => data_o <= x"00000004";
      when 592 => data_o <= x"FFFFF218";
      when 593 => data_o <= x"0000000A";
      when 594 => data_o <= x"0000A488";
      when 595 => data_o <= x"0000094C";
      when 596 => data_o <= x"FFFFF338";
      when 597 => data_o <= x"00000006";
      when 598 => data_o <= x"FFFFF22C";
      when 599 => data_o <= x"FFFFF334";
      when 600 => data_o <= x"00000538";
      when 601 => data_o <= x"00000001";
      when 602 => data_o <= x"0000000C";
      when 603 => data_o <= x"FFFFF26C";
      when 604 => data_o <= x"0000000C";
      when 605 => data_o <= x"00000001";
      when 606 => data_o <= x"FFFFF248";
      when 607 => data_o <= x"001A0001";
      when 608 => data_o <= x"00000003";
      when 609 => data_o <= x"FFFFF25C";
      when 610 => data_o <= x"0000A44C";
      when 611 => data_o <= x"00050003";
      when 612 => data_o <= x"FFFFF334";
      when 613 => data_o <= x"00000001";
      when 614 => data_o <= x"FFFFF334";
      when 615 => data_o <= x"0000A464";
      when 616 => data_o <= x"00000000";
      when 617 => data_o <= x"FFFFF338";
      when 618 => data_o <= x"F4000DFF";
      when 619 => data_o <= x"D01D0920";
      when 620 => data_o <= x"74000091";
      when 621 => data_o <= x"F4000928";
      when 622 => data_o <= x"9B9E4910";
      when 623 => data_o <= x"103F1FF0";
      when 624 => data_o <= x"28120000";
      when 625 => data_o <= x"E9500274";
      when 626 => data_o <= x"7E629D6F";
      when 627 => data_o <= x"5400026E";
      when 628 => data_o <= x"2BD00D97";
      when 629 => data_o <= x"D27EC800";
      when 630 => data_o <= x"F4000DFF";
      when 631 => data_o <= x"D3FF4EFF";
      when 632 => data_o <= x"D37F4E13";
      when 633 => data_o <= x"D2FF4D97";
      when 634 => data_o <= x"D2E7C800";
      when 635 => data_o <= x"F4010000";
      when 636 => data_o <= x"F4000DDF";
      when 637 => data_o <= x"D27EC800";
      when 638 => data_o <= x"F4018000";
      when 639 => data_o <= x"F4000DE3";
      when 640 => data_o <= x"D27EC220";
      when 641 => data_o <= x"7400026A";
      when 642 => data_o <= x"7400023B";
      when 643 => data_o <= x"54000108";
      when 644 => data_o <= x"7400026A";
      when 645 => data_o <= x"7400023B";
      when 646 => data_o <= x"54000108";
      when others => data_o <= x"00000000";
    end case;
  end if;
end process;

END ARCHITECTURE RTL;
