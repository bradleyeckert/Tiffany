library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

-- Single-port synchronous-read ROM

ENTITY ROM32 IS
generic (
  Size:  integer := 10                          -- log2 (cells)
);
port (
  clk:    in  std_logic;                        -- System clock
  addr:   in  std_logic_vector(Size-1 downto 0);
  data_o: out std_logic_vector(31 downto 0)     -- read data
);
END ROM32;

ARCHITECTURE RTL OF ROM32 IS
signal address: integer range 0 to 2**Size-1;
begin
address <= to_integer(unsigned(addr));

process (clk) begin
  if rising_edge(clk) then
    case address is
      when   0 => data_o <= x"54000A28";
      when   1 => data_o <= x"54000A2B";
      when   2 => data_o <= x"540001CE";
      when   3 => data_o <= x"85B693ED";
      when   4 => data_o <= x"000028B8";
      when   5 => data_o <= x"D090C220";
      when   6 => data_o <= x"9FB08800";
      when   7 => data_o <= x"3FB08800";
      when   8 => data_o <= x"5FB08800";
      when   9 => data_o <= x"05FB8328";
      when  10 => data_o <= x"9FB08800";
      when  11 => data_o <= x"05FD8328";
      when  12 => data_o <= x"3FB08800";
      when  13 => data_o <= x"D0908800";
      when  14 => data_o <= x"D09D0220";
      when  15 => data_o <= x"D21D0220";
      when  16 => data_o <= x"10408800";
      when  17 => data_o <= x"7FC2BC08";
      when  18 => data_o <= x"F1FF0A08";
      when  19 => data_o <= x"F3908800";
      when  20 => data_o <= x"F3B08800";
      when  21 => data_o <= x"F0AF1FF0";
      when  22 => data_o <= x"7DF08800";
      when  23 => data_o <= x"28AF0AF0";
      when  24 => data_o <= x"7FC08800";
      when  25 => data_o <= x"28A4BC7C";
      when  26 => data_o <= x"F12F1F08";
      when  27 => data_o <= x"EFB08800";
      when  28 => data_o <= x"E7908800";
      when  29 => data_o <= x"7FC2BC7C";
      when  30 => data_o <= x"7FC2BC2A";
      when  31 => data_o <= x"7DFE7928";
      when  32 => data_o <= x"2950001D";
      when  33 => data_o <= x"EFBEC220";
      when  34 => data_o <= x"07A08800";
      when  35 => data_o <= x"04220000";
      when  36 => data_o <= x"07005BD2";
      when  37 => data_o <= x"05B08800";
      when  38 => data_o <= x"90220000";
      when  39 => data_o <= x"6E408800";
      when  40 => data_o <= x"6E490220";
      when  41 => data_o <= x"92408800";
      when  42 => data_o <= x"D09B0220";
      when  43 => data_o <= x"24927D03";
      when  44 => data_o <= x"D1308800";
      when  45 => data_o <= x"9BCBBC08";
      when  46 => data_o <= x"9E7EC220";
      when  47 => data_o <= x"C3424800";
      when  48 => data_o <= x"08800000";
      when  49 => data_o <= x"D3CD13D2";
      when  50 => data_o <= x"7C220000";
      when  51 => data_o <= x"7DFF0A0C";
      when  52 => data_o <= x"F0A8C220";
      when  53 => data_o <= x"D1FD0928";
      when  54 => data_o <= x"E64C3B26";
      when  55 => data_o <= x"EC220000";
      when  56 => data_o <= x"C1500035";
      when  57 => data_o <= x"08800000";
      when  58 => data_o <= x"38220000";
      when  59 => data_o <= x"F4000004";
      when  60 => data_o <= x"66E08800";
      when  61 => data_o <= x"F4000008";
      when  62 => data_o <= x"66E08800";
      when  63 => data_o <= x"F400000C";
      when  64 => data_o <= x"A6EF4008";
      when  65 => data_o <= x"67424350";
      when  66 => data_o <= x"50220000";
      when  67 => data_o <= x"044119B8";
      when  68 => data_o <= x"F3B08800";
      when  69 => data_o <= x"F400000A";
      when  70 => data_o <= x"F4000DE7";
      when  71 => data_o <= x"D27EC220";
      when  72 => data_o <= x"F4000010";
      when  73 => data_o <= x"F4000DE7";
      when  74 => data_o <= x"D27EC220";
      when  75 => data_o <= x"B8800000";
      when  76 => data_o <= x"F4FFFFFF";
      when  77 => data_o <= x"4C220000";
      when  78 => data_o <= x"E79D0320";
      when  79 => data_o <= x"C3BEFB08";
      when  80 => data_o <= x"EFCD0928";
      when  81 => data_o <= x"87C7FC7C";
      when  82 => data_o <= x"7C220000";
      when  83 => data_o <= x"28A24AE4";
      when  84 => data_o <= x"E4320000";
      when  85 => data_o <= x"C3B7DF7E";
      when  86 => data_o <= x"EFBEE17E";
      when  87 => data_o <= x"2BC2B90C";
      when  88 => data_o <= x"4B90FC7C";
      when  89 => data_o <= x"F2C6C800";
      when  90 => data_o <= x"C3B7C220";
      when  91 => data_o <= x"ECAECAEC";
      when  92 => data_o <= x"85F08800";
      when  93 => data_o <= x"F400000C";
      when  94 => data_o <= x"46E08800";
      when  95 => data_o <= x"28AECAEC";
      when  96 => data_o <= x"7C220000";
      when  97 => data_o <= x"E796E420";
      when  98 => data_o <= x"EBB08800";
      when  99 => data_o <= x"EFB2A17E";
      when 100 => data_o <= x"28AD09D0";
      when 101 => data_o <= x"C3B7C220";
      when 102 => data_o <= x"7E17C220";
      when 103 => data_o <= x"281383F7";
      when 104 => data_o <= x"05F0CAD0";
      when 105 => data_o <= x"4DF08800";
      when 106 => data_o <= x"D090CCF5";
      when 107 => data_o <= x"4F427408";
      when 108 => data_o <= x"F150006A";
      when 109 => data_o <= x"E796EC20";
      when 110 => data_o <= x"EB4243B2";
      when 111 => data_o <= x"EEC08800";
      when 112 => data_o <= x"F150006D";
      when 113 => data_o <= x"D09D0800";
      when 114 => data_o <= x"C1500076";
      when 115 => data_o <= x"D09F1FF0";
      when 116 => data_o <= x"98A9DFA0";
      when 117 => data_o <= x"2BBEFB08";
      when 118 => data_o <= x"EFBEC220";
      when 119 => data_o <= x"D09D0800";
      when 120 => data_o <= x"C150007C";
      when 121 => data_o <= x"D09F1FF0";
      when 122 => data_o <= x"38A3DFA0";
      when 123 => data_o <= x"2BBEFB08";
      when 124 => data_o <= x"EFBEC220";
      when 125 => data_o <= x"D09D0800";
      when 126 => data_o <= x"C1500086";
      when 127 => data_o <= x"2417C3F0";
      when 128 => data_o <= x"483F0AD0";
      when 129 => data_o <= x"24800000";
      when 130 => data_o <= x"7F4274F0";
      when 131 => data_o <= x"D09D3CE4";
      when 132 => data_o <= x"DB93FB28";
      when 133 => data_o <= x"27054082";
      when 134 => data_o <= x"EFBEC220";
      when 135 => data_o <= x"7F9E5D6A";
      when 136 => data_o <= x"E950008B";
      when 137 => data_o <= x"29D0007D";
      when 138 => data_o <= x"5400008C";
      when 139 => data_o <= x"29D00077";
      when 140 => data_o <= x"08800000";
      when 141 => data_o <= x"E7A54092";
      when 142 => data_o <= x"F34249F0";
      when 143 => data_o <= x"7FC20000";
      when 144 => data_o <= x"4BC3E800";
      when 145 => data_o <= x"2BBEFB08";
      when 146 => data_o <= x"EFBEC220";
      when 147 => data_o <= x"07AEFB08";
      when 148 => data_o <= x"E7974031";
      when 149 => data_o <= x"F4000003";
      when 150 => data_o <= x"4FA54099";
      when 151 => data_o <= x"F4000000";
      when 152 => data_o <= x"5400008D";
      when 153 => data_o <= x"0416DF50";
      when 154 => data_o <= x"534249F0";
      when 155 => data_o <= x"4BC9E800";
      when 156 => data_o <= x"2BBEFB08";
      when 157 => data_o <= x"D09D30EE";
      when 158 => data_o <= x"F400003F";
      when 159 => data_o <= x"4F427C20";
      when 160 => data_o <= x"12803CEE";
      when 161 => data_o <= x"08800000";
      when 162 => data_o <= x"D09D30EE";
      when 163 => data_o <= x"F400003F";
      when 164 => data_o <= x"4F427C20";
      when 165 => data_o <= x"72803CEE";
      when 166 => data_o <= x"08800000";
      when 167 => data_o <= x"34000005";
      when 168 => data_o <= x"F0D00003";
      when 169 => data_o <= x"08800000";
      when 170 => data_o <= x"34000005";
      when 171 => data_o <= x"F3B08800";
      when 172 => data_o <= x"34000003";
      when 173 => data_o <= x"ECD00004";
      when 174 => data_o <= x"F0D00003";
      when 175 => data_o <= x"F0220000";
      when 176 => data_o <= x"E796DFE4";
      when 177 => data_o <= x"7DD0002F";
      when 178 => data_o <= x"7DD00038";
      when 179 => data_o <= x"29D000AC";
      when 180 => data_o <= x"F0AB0800";
      when 181 => data_o <= x"E95000B7";
      when 182 => data_o <= x"D0920000";
      when 183 => data_o <= x"F0AB0800";
      when 184 => data_o <= x"E95000BA";
      when 185 => data_o <= x"D0920000";
      when 186 => data_o <= x"08800000";
      when 187 => data_o <= x"05FE796C";
      when 188 => data_o <= x"7C17DD2F";
      when 189 => data_o <= x"7DD00038";
      when 190 => data_o <= x"29D000AC";
      when 191 => data_o <= x"F0AB0800";
      when 192 => data_o <= x"E95000C2";
      when 193 => data_o <= x"D0920000";
      when 194 => data_o <= x"F0AB0800";
      when 195 => data_o <= x"E95000C9";
      when 196 => data_o <= x"D09E4800";
      when 197 => data_o <= x"E95000C9";
      when 198 => data_o <= x"49FF0AF0";
      when 199 => data_o <= x"D090FCD0";
      when 200 => data_o <= x"27420000";
      when 201 => data_o <= x"2BB08800";
      when 202 => data_o <= x"06C05F20";
      when 203 => data_o <= x"E95000CE";
      when 204 => data_o <= x"D097DD35";
      when 205 => data_o <= x"28800000";
      when 206 => data_o <= x"7C1B0800";
      when 207 => data_o <= x"E95000D1";
      when 208 => data_o <= x"48320000";
      when 209 => data_o <= x"29D000AC";
      when 210 => data_o <= x"2BA540D4";
      when 211 => data_o <= x"F3427C20";
      when 212 => data_o <= x"08800000";
      when 213 => data_o <= x"E6CF15CA";
      when 214 => data_o <= x"740000D5";
      when 215 => data_o <= x"EC220000";
      when 216 => data_o <= x"740000D5";
      when 217 => data_o <= x"F3B08800";
      when 218 => data_o <= x"E797406D";
      when 219 => data_o <= x"EBC20000";
      when 220 => data_o <= x"EC220000";
      when 221 => data_o <= x"E79F1D6D";
      when 222 => data_o <= x"EBC20000";
      when 223 => data_o <= x"EC220000";
      when 224 => data_o <= x"E797406A";
      when 225 => data_o <= x"EBC20000";
      when 226 => data_o <= x"EC220000";
      when 227 => data_o <= x"E79F1D6A";
      when 228 => data_o <= x"EBC20000";
      when 229 => data_o <= x"EC220000";
      when 230 => data_o <= x"7FC483F0";
      when 231 => data_o <= x"2B424308";
      when 232 => data_o <= x"E742437C";
      when 233 => data_o <= x"D090CA20";
      when 234 => data_o <= x"5400006A";
      when 235 => data_o <= x"E796EC7C";
      when 236 => data_o <= x"7400002F";
      when 237 => data_o <= x"F1D0002F";
      when 238 => data_o <= x"740000A7";
      when 239 => data_o <= x"2BA540F1";
      when 240 => data_o <= x"74000035";
      when 241 => data_o <= x"08800000";
      when 242 => data_o <= x"7DD000EB";
      when 243 => data_o <= x"295000CA";
      when 244 => data_o <= x"740000F2";
      when 245 => data_o <= x"F3B08800";
      when 246 => data_o <= x"34000001";
      when 247 => data_o <= x"540000F7";
      when 248 => data_o <= x"08800000";
      when 249 => data_o <= x"F3D00000";
      when 250 => data_o <= x"D1F20000";
      when 251 => data_o <= x"E7A54105";
      when 252 => data_o <= x"F34274F0";
      when 253 => data_o <= x"38A6FD07";
      when 254 => data_o <= x"D0800000";
      when 255 => data_o <= x"25F07D01";
      when 256 => data_o <= x"4F427DED";
      when 257 => data_o <= x"94B88320";
      when 258 => data_o <= x"4FC71B28";
      when 259 => data_o <= x"C15000FF";
      when 260 => data_o <= x"EDF540FB";
      when 261 => data_o <= x"EFB2B408";
      when 262 => data_o <= x"E5FF4004";
      when 263 => data_o <= x"65FF4DEB";
      when 264 => data_o <= x"D2E7FD00";
      when 265 => data_o <= x"47D00DEB";
      when 266 => data_o <= x"D27EDD32";
      when 267 => data_o <= x"2BD00DEB";
      when 268 => data_o <= x"D27ECAEC";
      when 269 => data_o <= x"2816C220";
      when 270 => data_o <= x"07AEC220";
      when 271 => data_o <= x"F4000DEB";
      when 272 => data_o <= x"D2EBCA20";
      when 273 => data_o <= x"F4000DEB";
      when 274 => data_o <= x"D27ECAF0";
      when 275 => data_o <= x"7F7EFCEC";
      when 276 => data_o <= x"28AF0220";
      when 277 => data_o <= x"08800000";
      when 278 => data_o <= x"04D00002";
      when 279 => data_o <= x"08800000";
      when 280 => data_o <= x"F4000021";
      when 281 => data_o <= x"740000AA";
      when 282 => data_o <= x"74000116";
      when 283 => data_o <= x"0C800000";
      when 284 => data_o <= x"74000115";
      when 285 => data_o <= x"05D00116";
      when 286 => data_o <= x"7400006D";
      when 287 => data_o <= x"E950011C";
      when 288 => data_o <= x"EC220000";
      when 289 => data_o <= x"F3D0FFFF";
      when 290 => data_o <= x"4C334000";
      when 291 => data_o <= x"08800000";
      when 292 => data_o <= x"74000121";
      when 293 => data_o <= x"EC220000";
      when 294 => data_o <= x"74000115";
      when 295 => data_o <= x"F4060000";
      when 296 => data_o <= x"34000000";
      when 297 => data_o <= x"E9500126";
      when 298 => data_o <= x"F4010000";
      when 299 => data_o <= x"54000124";
      when 300 => data_o <= x"54000150";
      when 301 => data_o <= x"3950012C";
      when 302 => data_o <= x"040A0D02";
      when 303 => data_o <= x"4A325B1B";
      when 304 => data_o <= x"F40004B8";
      when 305 => data_o <= x"5400012D";
      when 306 => data_o <= x"F40004BB";
      when 307 => data_o <= x"5400012D";
      when 308 => data_o <= x"F4000000";
      when 309 => data_o <= x"34000000";
      when 310 => data_o <= x"54000115";
      when 311 => data_o <= x"74000134";
      when 312 => data_o <= x"E9500137";
      when 313 => data_o <= x"F4020000";
      when 314 => data_o <= x"34000000";
      when 315 => data_o <= x"08800000";
      when 316 => data_o <= x"00000498";
      when 317 => data_o <= x"000004C0";
      when 318 => data_o <= x"000004C8";
      when 319 => data_o <= x"000004D0";
      when 320 => data_o <= x"000004DC";
      when 321 => data_o <= x"F40004F0";
      when 322 => data_o <= x"F4000DCF";
      when 323 => data_o <= x"D27EC220";
      when 324 => data_o <= x"104F4DCF";
      when 325 => data_o <= x"D2E0EE7E";
      when 326 => data_o <= x"F4000000";
      when 327 => data_o <= x"54000144";
      when 328 => data_o <= x"F4000001";
      when 329 => data_o <= x"54000144";
      when 330 => data_o <= x"F4000002";
      when 331 => data_o <= x"54000144";
      when 332 => data_o <= x"F4000003";
      when 333 => data_o <= x"54000144";
      when 334 => data_o <= x"F4000004";
      when 335 => data_o <= x"54000144";
      when 336 => data_o <= x"07AEFB08";
      when 337 => data_o <= x"D0920000";
      when 338 => data_o <= x"25F38800";
      when 339 => data_o <= x"74000146";
      when 340 => data_o <= x"2B054152";
      when 341 => data_o <= x"EFB08800";
      when 342 => data_o <= x"F4000020";
      when 343 => data_o <= x"54000146";
      when 344 => data_o <= x"C3B08800";
      when 345 => data_o <= x"74000156";
      when 346 => data_o <= x"D09D0800";
      when 347 => data_o <= x"54000158";
      when 348 => data_o <= x"08800000";
      when 349 => data_o <= x"07D00009";
      when 350 => data_o <= x"D03B3D06";
      when 351 => data_o <= x"D130FD37";
      when 352 => data_o <= x"0C220000";
      when 353 => data_o <= x"F4000CCB";
      when 354 => data_o <= x"D3D00D97";
      when 355 => data_o <= x"D27EC220";
      when 356 => data_o <= x"F4000D97";
      when 357 => data_o <= x"D017EED0";
      when 358 => data_o <= x"27404A9C";
      when 359 => data_o <= x"ECFEC220";
      when 360 => data_o <= x"07D00DE7";
      when 361 => data_o <= x"D2E7C800";
      when 362 => data_o <= x"E9500171";
      when 363 => data_o <= x"F4000000";
      when 364 => data_o <= x"49D000AC";
      when 365 => data_o <= x"2BC7DDAC";
      when 366 => data_o <= x"F1D0015D";
      when 367 => data_o <= x"74000164";
      when 368 => data_o <= x"28220000";
      when 369 => data_o <= x"29D000AC";
      when 370 => data_o <= x"F1D0015D";
      when 371 => data_o <= x"74000164";
      when 372 => data_o <= x"0416C220";
      when 373 => data_o <= x"74000168";
      when 374 => data_o <= x"E7974031";
      when 375 => data_o <= x"93A54175";
      when 376 => data_o <= x"08800000";
      when 377 => data_o <= x"B3A5417C";
      when 378 => data_o <= x"F400002D";
      when 379 => data_o <= x"74000164";
      when 380 => data_o <= x"08800000";
      when 381 => data_o <= x"EFBF4D97";
      when 382 => data_o <= x"D2EF4CCB";
      when 383 => data_o <= x"D39D090E";
      when 384 => data_o <= x"E7424320";
      when 385 => data_o <= x"74000158";
      when 386 => data_o <= x"5400012C";
      when 387 => data_o <= x"7C17DD38";
      when 388 => data_o <= x"74000161";
      when 389 => data_o <= x"74000175";
      when 390 => data_o <= x"29D00179";
      when 391 => data_o <= x"7400017D";
      when 392 => data_o <= x"29500180";
      when 393 => data_o <= x"F4000000";
      when 394 => data_o <= x"F1500183";
      when 395 => data_o <= x"7DD00024";
      when 396 => data_o <= x"29500183";
      when 397 => data_o <= x"F4000000";
      when 398 => data_o <= x"74000183";
      when 399 => data_o <= x"54000156";
      when 400 => data_o <= x"F4000000";
      when 401 => data_o <= x"5400018D";
      when 402 => data_o <= x"F4000DE7";
      when 403 => data_o <= x"D2EF400A";
      when 404 => data_o <= x"6FA54196";
      when 405 => data_o <= x"54000190";
      when 406 => data_o <= x"74000024";
      when 407 => data_o <= x"5400018D";
      when 408 => data_o <= x"B9500192";
      when 409 => data_o <= x"74000161";
      when 410 => data_o <= x"D0920000";
      when 411 => data_o <= x"7DD00168";
      when 412 => data_o <= x"28920000";
      when 413 => data_o <= x"C150019B";
      when 414 => data_o <= x"EDD00175";
      when 415 => data_o <= x"5400017D";
      when 416 => data_o <= x"F4000DE7";
      when 417 => data_o <= x"D2E7DD48";
      when 418 => data_o <= x"F4000000";
      when 419 => data_o <= x"F1D00199";
      when 420 => data_o <= x"2BD00DE7";
      when 421 => data_o <= x"D27EC800";
      when 422 => data_o <= x"7400012C";
      when 423 => data_o <= x"54000156";
      when 424 => data_o <= x"7C104A0C";
      when 425 => data_o <= x"7C800000";
      when 426 => data_o <= x"0526C800";
      when 427 => data_o <= x"E95001CC";
      when 428 => data_o <= x"74000115";
      when 429 => data_o <= x"7400014C";
      when 430 => data_o <= x"E95001AC";
      when 431 => data_o <= x"7400014E";
      when 432 => data_o <= x"07D0000D";
      when 433 => data_o <= x"6E420000";
      when 434 => data_o <= x"E95001B5";
      when 435 => data_o <= x"ECAEFCD0";
      when 436 => data_o <= x"24308800";
      when 437 => data_o <= x"07D00008";
      when 438 => data_o <= x"6E420000";
      when 439 => data_o <= x"E95001C1";
      when 440 => data_o <= x"EF9E5B20";
      when 441 => data_o <= x"E95001C0";
      when 442 => data_o <= x"D09D0800";
      when 443 => data_o <= x"540001BE";
      when 444 => data_o <= x"445B1B07";
      when 445 => data_o <= x"445B1B20";
      when 446 => data_o <= x"F40006F0";
      when 447 => data_o <= x"39D0012C";
      when 448 => data_o <= x"540001CB";
      when 449 => data_o <= x"07D00020";
      when 450 => data_o <= x"D090C800";
      when 451 => data_o <= x"C15001CA";
      when 452 => data_o <= x"EFD00DB1";
      when 453 => data_o <= x"D3690800";
      when 454 => data_o <= x"E95001C8";
      when 455 => data_o <= x"05D00146";
      when 456 => data_o <= x"F0F20000";
      when 457 => data_o <= x"540001CB";
      when 458 => data_o <= x"EFB20000";
      when 459 => data_o <= x"540001AA";
      when 460 => data_o <= x"2BBF3427";
      when 461 => data_o <= x"08800000";
      when 462 => data_o <= x"0715410E";
      when 463 => data_o <= x"F4080000";
      when 464 => data_o <= x"34000000";
      when 465 => data_o <= x"93A541CF";
      when 466 => data_o <= x"F4030000";
      when 467 => data_o <= x"54000121";
      when 468 => data_o <= x"F4000D97";
      when 469 => data_o <= x"D01B9FF0";
      when 470 => data_o <= x"7DF741CF";
      when 471 => data_o <= x"ED29FB28";
      when 472 => data_o <= x"39F39FD8";
      when 473 => data_o <= x"740001CF";
      when 474 => data_o <= x"ECA741CF";
      when 475 => data_o <= x"ECA28320";
      when 476 => data_o <= x"740001CF";
      when 477 => data_o <= x"ECAF4D97";
      when 478 => data_o <= x"D27EC220";
      when 479 => data_o <= x"F4000005";
      when 480 => data_o <= x"740001CF";
      when 481 => data_o <= x"EFD001FF";
      when 482 => data_o <= x"540001CF";
      when 483 => data_o <= x"740001DF";
      when 484 => data_o <= x"F4000001";
      when 485 => data_o <= x"4E420000";
      when 486 => data_o <= x"E95001E3";
      when 487 => data_o <= x"08800000";
      when 488 => data_o <= x"F400009F";
      when 489 => data_o <= x"740001CF";
      when 490 => data_o <= x"05B741CF";
      when 491 => data_o <= x"05B741CF";
      when 492 => data_o <= x"05B541CF";
      when 493 => data_o <= x"F4000106";
      when 494 => data_o <= x"740001CF";
      when 495 => data_o <= x"EFD00020";
      when 496 => data_o <= x"F4000100";
      when 497 => data_o <= x"740001D4";
      when 498 => data_o <= x"F4000104";
      when 499 => data_o <= x"740001CF";
      when 500 => data_o <= x"ED5001E3";
      when 501 => data_o <= x"F40000FF";
      when 502 => data_o <= x"740001CF";
      when 503 => data_o <= x"F0F08800";
      when 504 => data_o <= x"F4000106";
      when 505 => data_o <= x"740001CF";
      when 506 => data_o <= x"EFCF4002";
      when 507 => data_o <= x"F4000000";
      when 508 => data_o <= x"740001D4";
      when 509 => data_o <= x"D09D1F38";
      when 510 => data_o <= x"4A420000";
      when 511 => data_o <= x"E9500206";
      when 512 => data_o <= x"F4000100";
      when 513 => data_o <= x"0DD001CF";
      when 514 => data_o <= x"EFD00104";
      when 515 => data_o <= x"740001CF";
      when 516 => data_o <= x"EDD001E3";
      when 517 => data_o <= x"2BB08800";
      when 518 => data_o <= x"740001CF";
      when 519 => data_o <= x"ECA541FD";
      when 520 => data_o <= x"08800000";
      when 521 => data_o <= x"F4000D97";
      when 522 => data_o <= x"D2E7F920";
      when 523 => data_o <= x"F400000B";
      when 524 => data_o <= x"F4000000";
      when 525 => data_o <= x"05F741D4";
      when 526 => data_o <= x"29D001CF";
      when 527 => data_o <= x"EDD0003B";
      when 528 => data_o <= x"E7424800";
      when 529 => data_o <= x"7CEF4D97";
      when 530 => data_o <= x"D017C800";
      when 531 => data_o <= x"740001F5";
      when 532 => data_o <= x"ECAD9D31";
      when 533 => data_o <= x"F40000FF";
      when 534 => data_o <= x"6FA54219";
      when 535 => data_o <= x"F400003B";
      when 536 => data_o <= x"D1D0010E";
      when 537 => data_o <= x"28920000";
      when 538 => data_o <= x"C1500211";
      when 539 => data_o <= x"EFBF41FF";
      when 540 => data_o <= x"740001CF";
      when 541 => data_o <= x"ECAF4D97";
      when 542 => data_o <= x"D27EC220";
      when 543 => data_o <= x"74000209";
      when 544 => data_o <= x"07AEFBEE";
      when 545 => data_o <= x"E74F40FF";
      when 546 => data_o <= x"4C9E5F20";
      when 547 => data_o <= x"740000DA";
      when 548 => data_o <= x"7FCE5220";
      when 549 => data_o <= x"740001F8";
      when 550 => data_o <= x"F120CA28";
      when 551 => data_o <= x"F3424320";
      when 552 => data_o <= x"54000220";
      when 553 => data_o <= x"08800000";
      when 554 => data_o <= x"F3D00D97";
      when 555 => data_o <= x"D27EC800";
      when 556 => data_o <= x"F4000D97";
      when 557 => data_o <= x"D3CF4004";
      when 558 => data_o <= x"5400021F";
      when 559 => data_o <= x"F400000B";
      when 560 => data_o <= x"F4000000";
      when 561 => data_o <= x"740001D4";
      when 562 => data_o <= x"05D001CF";
      when 563 => data_o <= x"EFD00D97";
      when 564 => data_o <= x"D1D001F5";
      when 565 => data_o <= x"740001F5";
      when 566 => data_o <= x"740001F5";
      when 567 => data_o <= x"740001F5";
      when 568 => data_o <= x"EFD001FF";
      when 569 => data_o <= x"740001CF";
      when 570 => data_o <= x"EFD00D97";
      when 571 => data_o <= x"D2E08800";
      when 572 => data_o <= x"07D08000";
      when 573 => data_o <= x"D090C800";
      when 574 => data_o <= x"C3B9FB08";
      when 575 => data_o <= x"ED50022A";
      when 576 => data_o <= x"07D08000";
      when 577 => data_o <= x"D090C800";
      when 578 => data_o <= x"C1500247";
      when 579 => data_o <= x"EFCF4D97";
      when 580 => data_o <= x"D017CFEC";
      when 581 => data_o <= x"2BCF4001";
      when 582 => data_o <= x"5400021F";
      when 583 => data_o <= x"EDFD3DFF";
      when 584 => data_o <= x"4D2F4003";
      when 585 => data_o <= x"4C410420";
      when 586 => data_o <= x"7400009D";
      when 587 => data_o <= x"D0AF4003";
      when 588 => data_o <= x"D139FB08";
      when 589 => data_o <= x"07D08000";
      when 590 => data_o <= x"D090C800";
      when 591 => data_o <= x"C1500251";
      when 592 => data_o <= x"ED50021F";
      when 593 => data_o <= x"EF424800";
      when 594 => data_o <= x"7F9DB920";
      when 595 => data_o <= x"74000240";
      when 596 => data_o <= x"27C27C28";
      when 597 => data_o <= x"27054252";
      when 598 => data_o <= x"EFBEC220";
      when 599 => data_o <= x"F4000000";
      when 600 => data_o <= x"F4000D9C";
      when 601 => data_o <= x"D0FEC220";
      when 602 => data_o <= x"F4000001";
      when 603 => data_o <= x"F4000D9C";
      when 604 => data_o <= x"D0FEC220";
      when 605 => data_o <= x"F4000D9C";
      when 606 => data_o <= x"D3620000";
      when 607 => data_o <= x"E9500262";
      when 608 => data_o <= x"F4000DDF";
      when 609 => data_o <= x"D0220000";
      when 610 => data_o <= x"F4000DDB";
      when 611 => data_o <= x"D0220000";
      when 612 => data_o <= x"05FB8800";
      when 613 => data_o <= x"7400023C";
      when 614 => data_o <= x"F4000004";
      when 615 => data_o <= x"29500009";
      when 616 => data_o <= x"F4000DDF";
      when 617 => data_o <= x"D1500264";
      when 618 => data_o <= x"F4000DE3";
      when 619 => data_o <= x"D1500264";
      when 620 => data_o <= x"F4000DDB";
      when 621 => data_o <= x"D017EE9C";
      when 622 => data_o <= x"EFD00004";
      when 623 => data_o <= x"29500009";
      when 624 => data_o <= x"F4000D9C";
      when 625 => data_o <= x"D3620000";
      when 626 => data_o <= x"E9500274";
      when 627 => data_o <= x"54000268";
      when 628 => data_o <= x"5400026C";
      when 629 => data_o <= x"05FB8800";
      when 630 => data_o <= x"74000240";
      when 631 => data_o <= x"4AE24A9C";
      when 632 => data_o <= x"EC220000";
      when 633 => data_o <= x"F4000DDF";
      when 634 => data_o <= x"D1500275";
      when 635 => data_o <= x"F4000DE3";
      when 636 => data_o <= x"D1500275";
      when 637 => data_o <= x"F4000DDB";
      when 638 => data_o <= x"D017EE3C";
      when 639 => data_o <= x"EFD00001";
      when 640 => data_o <= x"29500009";
      when 641 => data_o <= x"F4000D9C";
      when 642 => data_o <= x"D3620000";
      when 643 => data_o <= x"E9500285";
      when 644 => data_o <= x"54000279";
      when 645 => data_o <= x"5400027D";
      when 646 => data_o <= x"E7D00DDB";
      when 647 => data_o <= x"D2E6D308";
      when 648 => data_o <= x"F4000DDF";
      when 649 => data_o <= x"D2EF3D00";
      when 650 => data_o <= x"D1D00268";
      when 651 => data_o <= x"06E90800";
      when 652 => data_o <= x"74000286";
      when 653 => data_o <= x"E950028F";
      when 654 => data_o <= x"8550028B";
      when 655 => data_o <= x"04174268";
      when 656 => data_o <= x"06E92420";
      when 657 => data_o <= x"74000286";
      when 658 => data_o <= x"E9500295";
      when 659 => data_o <= x"99D00268";
      when 660 => data_o <= x"54000290";
      when 661 => data_o <= x"08800000";
      when 662 => data_o <= x"F4000DC7";
      when 663 => data_o <= x"D2EF4DBF";
      when 664 => data_o <= x"D27EC800";
      when 665 => data_o <= x"F4000D97";
      when 666 => data_o <= x"D3D000CC";
      when 667 => data_o <= x"74000093";
      when 668 => data_o <= x"F4000000";
      when 669 => data_o <= x"A4800000";
      when 670 => data_o <= x"74000288";
      when 671 => data_o <= x"7F42520C";
      when 672 => data_o <= x"514F39F0";
      when 673 => data_o <= x"7400023C";
      when 674 => data_o <= x"2BC90800";
      when 675 => data_o <= x"E950029E";
      when 676 => data_o <= x"EC220000";
      when 677 => data_o <= x"540002EC";
      when 678 => data_o <= x"540002F7";
      when 679 => data_o <= x"F4000000";
      when 680 => data_o <= x"F4000DA7";
      when 681 => data_o <= x"D27EFD1A";
      when 682 => data_o <= x"F4000DB5";
      when 683 => data_o <= x"D17EFD00";
      when 684 => data_o <= x"F4000DB6";
      when 685 => data_o <= x"D0FEC220";
      when 686 => data_o <= x"F3D00DB5";
      when 687 => data_o <= x"D367409D";
      when 688 => data_o <= x"F4000DA7";
      when 689 => data_o <= x"D2E0C320";
      when 690 => data_o <= x"F4000DA7";
      when 691 => data_o <= x"D27EC220";
      when 692 => data_o <= x"740002A5";
      when 693 => data_o <= x"F4000DB5";
      when 694 => data_o <= x"D3693920";
      when 695 => data_o <= x"F400003C";
      when 696 => data_o <= x"4D320000";
      when 697 => data_o <= x"E95002BB";
      when 698 => data_o <= x"740002A6";
      when 699 => data_o <= x"F4000000";
      when 700 => data_o <= x"740002AE";
      when 701 => data_o <= x"F4000DB5";
      when 702 => data_o <= x"D3604800";
      when 703 => data_o <= x"E95002C4";
      when 704 => data_o <= x"F4000006";
      when 705 => data_o <= x"D090C1B0";
      when 706 => data_o <= x"D13F4DB5";
      when 707 => data_o <= x"D0FEC220";
      when 708 => data_o <= x"ED5002A6";
      when 709 => data_o <= x"F1D002A5";
      when 710 => data_o <= x"F4000001";
      when 711 => data_o <= x"F4000DB5";
      when 712 => data_o <= x"D3605F20";
      when 713 => data_o <= x"7400009D";
      when 714 => data_o <= x"E5D0006D";
      when 715 => data_o <= x"2A474031";
      when 716 => data_o <= x"E95002CE";
      when 717 => data_o <= x"740002A6";
      when 718 => data_o <= x"740002AE";
      when 719 => data_o <= x"F4000DB5";
      when 720 => data_o <= x"D36F4018";
      when 721 => data_o <= x"7400009D";
      when 722 => data_o <= x"F4000DDF";
      when 723 => data_o <= x"D2E0C800";
      when 724 => data_o <= x"F4000DAF";
      when 725 => data_o <= x"D27EFD00";
      when 726 => data_o <= x"F4000DB5";
      when 727 => data_o <= x"D0FEC800";
      when 728 => data_o <= x"540002A6";
      when 729 => data_o <= x"05FC3424";
      when 730 => data_o <= x"F5FFFFFF";
      when 731 => data_o <= x"D04E5320";
      when 732 => data_o <= x"E95002E4";
      when 733 => data_o <= x"ECA07D18";
      when 734 => data_o <= x"740000A2";
      when 735 => data_o <= x"F400003D";
      when 736 => data_o <= x"740002C5";
      when 737 => data_o <= x"F4FFFFFF";
      when 738 => data_o <= x"4FD00025";
      when 739 => data_o <= x"540002C5";
      when 740 => data_o <= x"2AC20000";
      when 741 => data_o <= x"E95002EA";
      when 742 => data_o <= x"D09D3D3D";
      when 743 => data_o <= x"740002C5";
      when 744 => data_o <= x"F4000034";
      when 745 => data_o <= x"540002B4";
      when 746 => data_o <= x"F400003D";
      when 747 => data_o <= x"540002C5";
      when 748 => data_o <= x"F4000DB4";
      when 749 => data_o <= x"D3620000";
      when 750 => data_o <= x"E95002F4";
      when 751 => data_o <= x"F4000000";
      when 752 => data_o <= x"F4000DB4";
      when 753 => data_o <= x"D0FEC800";
      when 754 => data_o <= x"F4000DAB";
      when 755 => data_o <= x"D2E742D9";
      when 756 => data_o <= x"F4000000";
      when 757 => data_o <= x"F4000DB6";
      when 758 => data_o <= x"D0FEC220";
      when 759 => data_o <= x"740002A5";
      when 760 => data_o <= x"F4000DB5";
      when 761 => data_o <= x"D36F4015";
      when 762 => data_o <= x"E7424320";
      when 763 => data_o <= x"C3BEC220";
      when 764 => data_o <= x"EFA542FF";
      when 765 => data_o <= x"F4000008";
      when 766 => data_o <= x"740002B4";
      when 767 => data_o <= x"F4000DA7";
      when 768 => data_o <= x"D2E74268";
      when 769 => data_o <= x"540002A7";
      when 770 => data_o <= x"740002A5";
      when 771 => data_o <= x"F5FFFFFF";
      when 772 => data_o <= x"D04E5320";
      when 773 => data_o <= x"E9500307";
      when 774 => data_o <= x"540002D9";
      when 775 => data_o <= x"F4000DAB";
      when 776 => data_o <= x"D27EFD01";
      when 777 => data_o <= x"F4000DB4";
      when 778 => data_o <= x"D0FEC220";
      when 779 => data_o <= x"514F401D";
      when 780 => data_o <= x"740002C5";
      when 781 => data_o <= x"F4000DA3";
      when 782 => data_o <= x"D2EF4004";
      when 783 => data_o <= x"0F6F4080";
      when 784 => data_o <= x"4FD00DB6";
      when 785 => data_o <= x"D0FEC220";
      when 786 => data_o <= x"F4000DB6";
      when 787 => data_o <= x"D3620000";
      when 788 => data_o <= x"E9500320";
      when 789 => data_o <= x"F4000DAF";
      when 790 => data_o <= x"D1D0004B";
      when 791 => data_o <= x"F4000008";
      when 792 => data_o <= x"F4000DAC";
      when 793 => data_o <= x"D367409D";
      when 794 => data_o <= x"D3C7423C";
      when 795 => data_o <= x"F4000000";
      when 796 => data_o <= x"F4000DB6";
      when 797 => data_o <= x"D0FEFD00";
      when 798 => data_o <= x"F4000DAF";
      when 799 => data_o <= x"D27EC220";
      when 800 => data_o <= x"F4000002";
      when 801 => data_o <= x"540002B4";
      when 802 => data_o <= x"F4000DE7";
      when 803 => data_o <= x"D017EE20";
      when 804 => data_o <= x"F400003B";
      when 805 => data_o <= x"74000146";
      when 806 => data_o <= x"F1D00045";
      when 807 => data_o <= x"F4000000";
      when 808 => data_o <= x"7400018B";
      when 809 => data_o <= x"2A7EC220";
      when 810 => data_o <= x"F4000DB0";
      when 811 => data_o <= x"D36E8AEE";
      when 812 => data_o <= x"08800000";
      when 813 => data_o <= x"F4000000";
      when 814 => data_o <= x"F4000DB0";
      when 815 => data_o <= x"D0FEC220";
      when 816 => data_o <= x"F4000001";
      when 817 => data_o <= x"F4000DB0";
      when 818 => data_o <= x"D0FEC220";
      when 819 => data_o <= x"F400001B";
      when 820 => data_o <= x"74000146";
      when 821 => data_o <= x"F400005B";
      when 822 => data_o <= x"74000146";
      when 823 => data_o <= x"54000146";
      when 824 => data_o <= x"F4000030";
      when 825 => data_o <= x"54000333";
      when 826 => data_o <= x"F4000031";
      when 827 => data_o <= x"54000333";
      when 828 => data_o <= x"F400006D";
      when 829 => data_o <= x"54000146";
      when 830 => data_o <= x"7400032A";
      when 831 => data_o <= x"74000338";
      when 832 => data_o <= x"5400033C";
      when 833 => data_o <= x"7400033A";
      when 834 => data_o <= x"74000322";
      when 835 => data_o <= x"5400033C";
      when 836 => data_o <= x"74000338";
      when 837 => data_o <= x"74000322";
      when 838 => data_o <= x"5400033C";
      when 839 => data_o <= x"7400032A";
      when 840 => data_o <= x"F4000023";
      when 841 => data_o <= x"54000341";
      when 842 => data_o <= x"7400032A";
      when 843 => data_o <= x"F400001F";
      when 844 => data_o <= x"54000341";
      when 845 => data_o <= x"7400032A";
      when 846 => data_o <= x"F4000020";
      when 847 => data_o <= x"54000341";
      when 848 => data_o <= x"7400032A";
      when 849 => data_o <= x"F4000021";
      when 850 => data_o <= x"54000341";
      when 851 => data_o <= x"7400032A";
      when 852 => data_o <= x"F4000021";
      when 853 => data_o <= x"54000344";
      when 854 => data_o <= x"5400033E";
      when 855 => data_o <= x"28242D24";
      when 856 => data_o <= x"28202D20";
      when 857 => data_o <= x"2E212A21";
      when 858 => data_o <= x"28212C21";
      when 859 => data_o <= x"F4000DB0";
      when 860 => data_o <= x"D36EBB08";
      when 861 => data_o <= x"07D00001";
      when 862 => data_o <= x"4FA54362";
      when 863 => data_o <= x"EFD00028";
      when 864 => data_o <= x"F400001F";
      when 865 => data_o <= x"54000364";
      when 866 => data_o <= x"F4000D5C";
      when 867 => data_o <= x"0CEF36F0";
      when 868 => data_o <= x"7400033A";
      when 869 => data_o <= x"74000322";
      when 870 => data_o <= x"74000322";
      when 871 => data_o <= x"5400033C";
      when 872 => data_o <= x"7400003F";
      when 873 => data_o <= x"74000022";
      when 874 => data_o <= x"E9500370";
      when 875 => data_o <= x"D0920000";
      when 876 => data_o <= x"07425D43";
      when 877 => data_o <= x"74000192";
      when 878 => data_o <= x"2705436C";
      when 879 => data_o <= x"EC800000";
      when 880 => data_o <= x"54000372";
      when 881 => data_o <= x"70733C03";
      when 882 => data_o <= x"F4000DC4";
      when 883 => data_o <= x"39D0012C";
      when 884 => data_o <= x"54000148";
      when 885 => data_o <= x"F3D00003";
      when 886 => data_o <= x"D13F0800";
      when 887 => data_o <= x"07A5439A";
      when 888 => data_o <= x"E5D00347";
      when 889 => data_o <= x"F4000003";
      when 890 => data_o <= x"740001A0";
      when 891 => data_o <= x"74000350";
      when 892 => data_o <= x"E79F4004";
      when 893 => data_o <= x"05F740DA";
      when 894 => data_o <= x"2B9D090C";
      when 895 => data_o <= x"F4000009";
      when 896 => data_o <= x"740000AA";
      when 897 => data_o <= x"7C800000";
      when 898 => data_o <= x"07A54387";
      when 899 => data_o <= x"7E6F4007";
      when 900 => data_o <= x"740001A0";
      when 901 => data_o <= x"2B427420";
      when 902 => data_o <= x"54000382";
      when 903 => data_o <= x"EFB28800";
      when 904 => data_o <= x"74000158";
      when 905 => data_o <= x"E79F4010";
      when 906 => data_o <= x"740000DA";
      when 907 => data_o <= x"7400034D";
      when 908 => data_o <= x"07A54394";
      when 909 => data_o <= x"7CE07D20";
      when 910 => data_o <= x"F40000C0";
      when 911 => data_o <= x"740000E8";
      when 912 => data_o <= x"EBBF402E";
      when 913 => data_o <= x"74000146";
      when 914 => data_o <= x"2B427420";
      when 915 => data_o <= x"5400038C";
      when 916 => data_o <= x"EFBF4010";
      when 917 => data_o <= x"740000E6";
      when 918 => data_o <= x"F4000000";
      when 919 => data_o <= x"740000DD";
      when 920 => data_o <= x"74000148";
      when 921 => data_o <= x"54000377";
      when 922 => data_o <= x"EFB5433E";
      when 923 => data_o <= x"04800000";
      when 924 => data_o <= x"07A543A0";
      when 925 => data_o <= x"7FC2BC28";
      when 926 => data_o <= x"F1F7F424";
      when 927 => data_o <= x"D150039C";
      when 928 => data_o <= x"ECAF1F7E";
      when 929 => data_o <= x"28AF1F04";
      when 930 => data_o <= x"07A543A6";
      when 931 => data_o <= x"28AF1FF0";
      when 932 => data_o <= x"7FC2B424";
      when 933 => data_o <= x"D15003A2";
      when 934 => data_o <= x"EC220000";
      when 935 => data_o <= x"07D00061";
      when 936 => data_o <= x"F400007B";
      when 937 => data_o <= x"740000E8";
      when 938 => data_o <= x"F4000020";
      when 939 => data_o <= x"4F424308";
      when 940 => data_o <= x"7DD003A7";
      when 941 => data_o <= x"F4000030";
      when 942 => data_o <= x"D090C120";
      when 943 => data_o <= x"F400000A";
      when 944 => data_o <= x"F4000011";
      when 945 => data_o <= x"740000E8";
      when 946 => data_o <= x"91F07D09";
      when 947 => data_o <= x"74000070";
      when 948 => data_o <= x"F4000007";
      when 949 => data_o <= x"4F424328";
      when 950 => data_o <= x"E4A7406A";
      when 951 => data_o <= x"4C220000";
      when 952 => data_o <= x"07A543C6";
      when 953 => data_o <= x"7C17F620";
      when 954 => data_o <= x"F4000DE7";
      when 955 => data_o <= x"D2E743AC";
      when 956 => data_o <= x"E95003C5";
      when 957 => data_o <= x"F3D00DE7";
      when 958 => data_o <= x"D2E740A7";
      when 959 => data_o <= x"EDFF0AF0";
      when 960 => data_o <= x"F4000DE7";
      when 961 => data_o <= x"D2E740A7";
      when 962 => data_o <= x"74000033";
      when 963 => data_o <= x"2892B424";
      when 964 => data_o <= x"D15003B8";
      when 965 => data_o <= x"ECA28800";
      when 966 => data_o <= x"08800000";
      when 967 => data_o <= x"F4000DC7";
      when 968 => data_o <= x"D150002D";
      when 969 => data_o <= x"740003C7";
      when 970 => data_o <= x"F4000DBF";
      when 971 => data_o <= x"D2E540E6";
      when 972 => data_o <= x"7C800000";
      when 973 => data_o <= x"07A2BB08";
      when 974 => data_o <= x"E7649B90";
      when 975 => data_o <= x"E8AEC220";
      when 976 => data_o <= x"F4000001";
      when 977 => data_o <= x"740000E6";
      when 978 => data_o <= x"540003CD";
      when 979 => data_o <= x"08800000";
      when 980 => data_o <= x"7C800000";
      when 981 => data_o <= x"07A2BB08";
      when 982 => data_o <= x"E7649B20";
      when 983 => data_o <= x"E8AEC220";
      when 984 => data_o <= x"F4000001";
      when 985 => data_o <= x"740000E6";
      when 986 => data_o <= x"540003D5";
      when 987 => data_o <= x"08800000";
      when 988 => data_o <= x"740003C9";
      when 989 => data_o <= x"E5F7FC28";
      when 990 => data_o <= x"F1D003D4";
      when 991 => data_o <= x"29FF0AF0";
      when 992 => data_o <= x"E742437C";
      when 993 => data_o <= x"F0AF2490";
      when 994 => data_o <= x"F4000001";
      when 995 => data_o <= x"4F90C800";
      when 996 => data_o <= x"F4000DBF";
      when 997 => data_o <= x"D1500009";
      when 998 => data_o <= x"7DD003C9";
      when 999 => data_o <= x"E52F1F20";
      when 1000 => data_o <= x"740003CC";
      when 1001 => data_o <= x"ECAD090C";
      when 1002 => data_o <= x"F4000DBF";
      when 1003 => data_o <= x"D1D00009";
      when 1004 => data_o <= x"295003DC";
      when 1005 => data_o <= x"F4000020";
      when 1006 => data_o <= x"540003E6";
      when 1007 => data_o <= x"740003E6";
      when 1008 => data_o <= x"F4000D0B";
      when 1009 => data_o <= x"D017CFEC";
      when 1010 => data_o <= x"48E74077";
      when 1011 => data_o <= x"28220000";
      when 1012 => data_o <= x"F4000029";
      when 1013 => data_o <= x"740003DC";
      when 1014 => data_o <= x"5400012C";
      when 1015 => data_o <= x"740003ED";
      when 1016 => data_o <= x"EF608800";
      when 1017 => data_o <= x"7400003B";
      when 1018 => data_o <= x"E5B90800";
      when 1019 => data_o <= x"EBB05B08";
      when 1020 => data_o <= x"EF97DD3B";
      when 1021 => data_o <= x"7FCD0920";
      when 1022 => data_o <= x"7CE7FC38";
      when 1023 => data_o <= x"2BD00DB2";
      when 1024 => data_o <= x"D3690800";
      when 1025 => data_o <= x"E9500404";
      when 1026 => data_o <= x"740003A7";
      when 1027 => data_o <= x"F1D003A7";
      when 1028 => data_o <= x"6FA54407";
      when 1029 => data_o <= x"2BBEFB28";
      when 1030 => data_o <= x"28105B08";
      when 1031 => data_o <= x"28920000";
      when 1032 => data_o <= x"C15003FE";
      when 1033 => data_o <= x"EFBECAEC";
      when 1034 => data_o <= x"28908800";
      when 1035 => data_o <= x"BB9F401F";
      when 1036 => data_o <= x"7400006C";
      when 1037 => data_o <= x"F4000012";
      when 1038 => data_o <= x"D137410E";
      when 1039 => data_o <= x"E7A05B08";
      when 1040 => data_o <= x"05F84E20";
      when 1041 => data_o <= x"F400003F";
      when 1042 => data_o <= x"4DD003F9";
      when 1043 => data_o <= x"E9500415";
      when 1044 => data_o <= x"28220000";
      when 1045 => data_o <= x"29D0004B";
      when 1046 => data_o <= x"06420000";
      when 1047 => data_o <= x"E9500410";
      when 1048 => data_o <= x"08800000";
      when 1049 => data_o <= x"F4000DB7";
      when 1050 => data_o <= x"D3620000";
      when 1051 => data_o <= x"D09D0800";
      when 1052 => data_o <= x"C3BEC220";
      when 1053 => data_o <= x"7D210420";
      when 1054 => data_o <= x"F4000D9B";
      when 1055 => data_o <= x"D03B8800";
      when 1056 => data_o <= x"7400040B";
      when 1057 => data_o <= x"74000022";
      when 1058 => data_o <= x"E9500424";
      when 1059 => data_o <= x"2816FC08";
      when 1060 => data_o <= x"2815441B";
      when 1061 => data_o <= x"08800000";
      when 1062 => data_o <= x"F4000000";
      when 1063 => data_o <= x"F4000DB2";
      when 1064 => data_o <= x"D0FEC220";
      when 1065 => data_o <= x"F4000001";
      when 1066 => data_o <= x"F4000DB2";
      when 1067 => data_o <= x"D0FEC220";
      when 1068 => data_o <= x"740003ED";
      when 1069 => data_o <= x"74000419";
      when 1070 => data_o <= x"F2493D0C";
      when 1071 => data_o <= x"D135410E";
      when 1072 => data_o <= x"7400042C";
      when 1073 => data_o <= x"D21D154B";
      when 1074 => data_o <= x"E76F402D";
      when 1075 => data_o <= x"6E405F20";
      when 1076 => data_o <= x"E9500437";
      when 1077 => data_o <= x"F4000001";
      when 1078 => data_o <= x"740000E6";
      when 1079 => data_o <= x"28220000";
      when 1080 => data_o <= x"F4000000";
      when 1081 => data_o <= x"05D0001D";
      when 1082 => data_o <= x"740003B8";
      when 1083 => data_o <= x"924F400C";
      when 1084 => data_o <= x"D137410E";
      when 1085 => data_o <= x"EFB08800";
      when 1086 => data_o <= x"7FD00006";
      when 1087 => data_o <= x"7400009D";
      when 1088 => data_o <= x"28E07DC0";
      when 1089 => data_o <= x"4FD00080";
      when 1090 => data_o <= x"6E493D0C";
      when 1091 => data_o <= x"D137410E";
      when 1092 => data_o <= x"F400003F";
      when 1093 => data_o <= x"4FC7C32A";
      when 1094 => data_o <= x"E76F40F0";
      when 1095 => data_o <= x"7400006D";
      when 1096 => data_o <= x"E7D00001";
      when 1097 => data_o <= x"6E44C800";
      when 1098 => data_o <= x"E950044C";
      when 1099 => data_o <= x"EF608800";
      when 1100 => data_o <= x"E76F40E0";
      when 1101 => data_o <= x"7400006D";
      when 1102 => data_o <= x"E7D00002";
      when 1103 => data_o <= x"6E44C800";
      when 1104 => data_o <= x"E9500454";
      when 1105 => data_o <= x"ECEF401F";
      when 1106 => data_o <= x"4FC7443E";
      when 1107 => data_o <= x"EC220000";
      when 1108 => data_o <= x"E76F40F0";
      when 1109 => data_o <= x"7400006D";
      when 1110 => data_o <= x"E7D00003";
      when 1111 => data_o <= x"6E44C800";
      when 1112 => data_o <= x"E950045D";
      when 1113 => data_o <= x"ECEF401F";
      when 1114 => data_o <= x"4FC7443E";
      when 1115 => data_o <= x"7400043E";
      when 1116 => data_o <= x"EC220000";
      when 1117 => data_o <= x"F400000C";
      when 1118 => data_o <= x"D150010E";
      when 1119 => data_o <= x"74000432";
      when 1120 => data_o <= x"7F9E7D2E";
      when 1121 => data_o <= x"740003D4";
      when 1122 => data_o <= x"F3B20000";
      when 1123 => data_o <= x"E9500466";
      when 1124 => data_o <= x"F4000027";
      when 1125 => data_o <= x"D1D0010E";
      when 1126 => data_o <= x"07D00002";
      when 1127 => data_o <= x"74000070";
      when 1128 => data_o <= x"E9500483";
      when 1129 => data_o <= x"E79E43D0";
      when 1130 => data_o <= x"274DBCD8";
      when 1131 => data_o <= x"E5B93C20";
      when 1132 => data_o <= x"F4000027";
      when 1133 => data_o <= x"6E44C800";
      when 1134 => data_o <= x"E9500476";
      when 1135 => data_o <= x"F4000001";
      when 1136 => data_o <= x"740000E6";
      when 1137 => data_o <= x"D09D0800";
      when 1138 => data_o <= x"74000446";
      when 1139 => data_o <= x"2BA54475";
      when 1140 => data_o <= x"D0920000";
      when 1141 => data_o <= x"08800000";
      when 1142 => data_o <= x"E76F4024";
      when 1143 => data_o <= x"6E420000";
      when 1144 => data_o <= x"E9500483";
      when 1145 => data_o <= x"F4000DE7";
      when 1146 => data_o <= x"D2E7DD48";
      when 1147 => data_o <= x"F4000001";
      when 1148 => data_o <= x"740000E6";
      when 1149 => data_o <= x"74000438";
      when 1150 => data_o <= x"2BD00DE7";
      when 1151 => data_o <= x"D27ECA20";
      when 1152 => data_o <= x"E9500482";
      when 1153 => data_o <= x"D0920000";
      when 1154 => data_o <= x"08800000";
      when 1155 => data_o <= x"74000438";
      when 1156 => data_o <= x"2BA54486";
      when 1157 => data_o <= x"D0920000";
      when 1158 => data_o <= x"08800000";
      when 1159 => data_o <= x"740003ED";
      when 1160 => data_o <= x"07A544A2";
      when 1161 => data_o <= x"74000419";
      when 1162 => data_o <= x"E7A54491";
      when 1163 => data_o <= x"7400045F";
      when 1164 => data_o <= x"F4000DD7";
      when 1165 => data_o <= x"D2E20000";
      when 1166 => data_o <= x"E9500490";
      when 1167 => data_o <= x"74000302";
      when 1168 => data_o <= x"5400049E";
      when 1169 => data_o <= x"F3B04800";
      when 1170 => data_o <= x"F4000DA3";
      when 1171 => data_o <= x"D27EC800";
      when 1172 => data_o <= x"F4000DD7";
      when 1173 => data_o <= x"D2E92420";
      when 1174 => data_o <= x"F4000004";
      when 1175 => data_o <= x"4E1D090C";
      when 1176 => data_o <= x"7400004B";
      when 1177 => data_o <= x"04800000";
      when 1178 => data_o <= x"F4800000";
      when 1179 => data_o <= x"4E493D14";
      when 1180 => data_o <= x"D137410E";
      when 1181 => data_o <= x"74000032";
      when 1182 => data_o <= x"7400003F";
      when 1183 => data_o <= x"B3D00003";
      when 1184 => data_o <= x"D137410E";
      when 1185 => data_o <= x"54000487";
      when 1186 => data_o <= x"EFB08800";
      when 1187 => data_o <= x"F4000DA3";
      when 1188 => data_o <= x"D2ED21D0";
      when 1189 => data_o <= x"5400004B";
      when 1190 => data_o <= x"FFFFFFFF";
      when 1191 => data_o <= x"FFFFFFFF";
      when 1192 => data_o <= x"FFFFFFFF";
      when 1193 => data_o <= x"540004B3";
      when 1194 => data_o <= x"540004E7";
      when 1195 => data_o <= x"540004FA";
      when 1196 => data_o <= x"540004B5";
      when 1197 => data_o <= x"540004FE";
      when 1198 => data_o <= x"540004B0";
      when 1199 => data_o <= x"540004FC";
      when 1200 => data_o <= x"F4000DA3";
      when 1201 => data_o <= x"D2EF4010";
      when 1202 => data_o <= x"D090EE08";
      when 1203 => data_o <= x"740004A3";
      when 1204 => data_o <= x"54000032";
      when 1205 => data_o <= x"F4000DA3";
      when 1206 => data_o <= x"D2EF4014";
      when 1207 => data_o <= x"D090DD2D";
      when 1208 => data_o <= x"54000032";
      when 1209 => data_o <= x"F400000D";
      when 1210 => data_o <= x"D150010E";
      when 1211 => data_o <= x"740004AE";
      when 1212 => data_o <= x"A4220000";
      when 1213 => data_o <= x"04220000";
      when 1214 => data_o <= x"0C220000";
      when 1215 => data_o <= x"D090C220";
      when 1216 => data_o <= x"8C220000";
      when 1217 => data_o <= x"48220000";
      when 1218 => data_o <= x"4C220000";
      when 1219 => data_o <= x"E4220000";
      when 1220 => data_o <= x"28220000";
      when 1221 => data_o <= x"6C220000";
      when 1222 => data_o <= x"10220000";
      when 1223 => data_o <= x"30220000";
      when 1224 => data_o <= x"3C220000";
      when 1225 => data_o <= x"38220000";
      when 1226 => data_o <= x"38220000";
      when 1227 => data_o <= x"D8220000";
      when 1228 => data_o <= x"5C220000";
      when 1229 => data_o <= x"58220000";
      when 1230 => data_o <= x"78220000";
      when 1231 => data_o <= x"9C220000";
      when 1232 => data_o <= x"98220000";
      when 1233 => data_o <= x"B8220000";
      when 1234 => data_o <= x"70220000";
      when 1235 => data_o <= x"80220000";
      when 1236 => data_o <= x"A0220000";
      when 1237 => data_o <= x"50220000";
      when 1238 => data_o <= x"64220000";
      when 1239 => data_o <= x"D0220000";
      when 1240 => data_o <= x"BC220000";
      when 1241 => data_o <= x"44220000";
      when 1242 => data_o <= x"C4220000";
      when 1243 => data_o <= x"DC220000";
      when 1244 => data_o <= x"A4220000";
      when 1245 => data_o <= x"FC220000";
      when 1246 => data_o <= x"EC220000";
      when 1247 => data_o <= x"24220000";
      when 1248 => data_o <= x"24220000";
      when 1249 => data_o <= x"84220000";
      when 1250 => data_o <= x"7C220000";
      when 1251 => data_o <= x"F0220000";
      when 1252 => data_o <= x"90220000";
      when 1253 => data_o <= x"B0220000";
      when 1254 => data_o <= x"08800000";
      when 1255 => data_o <= x"740004A3";
      when 1256 => data_o <= x"9BD0001A";
      when 1257 => data_o <= x"06C20000";
      when 1258 => data_o <= x"E95004EF";
      when 1259 => data_o <= x"EFD00003";
      when 1260 => data_o <= x"4DF9BD1A";
      when 1261 => data_o <= x"28800000";
      when 1262 => data_o <= x"540004F3";
      when 1263 => data_o <= x"E79740A2";
      when 1264 => data_o <= x"F400003F";
      when 1265 => data_o <= x"4DFF4006";
      when 1266 => data_o <= x"D090CA20";
      when 1267 => data_o <= x"07D00002";
      when 1268 => data_o <= x"6E420000";
      when 1269 => data_o <= x"E95004F7";
      when 1270 => data_o <= x"EFBEFB08";
      when 1271 => data_o <= x"740002B4";
      when 1272 => data_o <= x"540004E9";
      when 1273 => data_o <= x"08800000";
      when 1274 => data_o <= x"740004A3";
      when 1275 => data_o <= x"5400030B";
      when 1276 => data_o <= x"740004AE";
      when 1277 => data_o <= x"54000302";
      when 1278 => data_o <= x"F4000DA3";
      when 1279 => data_o <= x"D2EF4014";
      when 1280 => data_o <= x"D090E620";
      when 1281 => data_o <= x"74000302";
      when 1282 => data_o <= x"B950030B";
      when 1283 => data_o <= x"740004AE";
      when 1284 => data_o <= x"540002B4";
      when 1285 => data_o <= x"F4000DB4";
      when 1286 => data_o <= x"D01D8800";
      when 1287 => data_o <= x"E950050E";
      when 1288 => data_o <= x"F4000000";
      when 1289 => data_o <= x"F0FEC800";
      when 1290 => data_o <= x"740004AE";
      when 1291 => data_o <= x"F4000DAB";
      when 1292 => data_o <= x"D2EF0800";
      when 1293 => data_o <= x"540002C5";
      when 1294 => data_o <= x"F400003A";
      when 1295 => data_o <= x"D150010E";
      when 1296 => data_o <= x"740002A5";
      when 1297 => data_o <= x"F4000DB5";
      when 1298 => data_o <= x"D3D00008";
      when 1299 => data_o <= x"7400006D";
      when 1300 => data_o <= x"E9500516";
      when 1301 => data_o <= x"740002A6";
      when 1302 => data_o <= x"740004AE";
      when 1303 => data_o <= x"540002B4";
      when 1304 => data_o <= x"740002A6";
      when 1305 => data_o <= x"740004AE";
      when 1306 => data_o <= x"540002B4";
      when 1307 => data_o <= x"740002A5";
      when 1308 => data_o <= x"540002A6";
      when 1309 => data_o <= x"740004AE";
      when 1310 => data_o <= x"74000302";
      when 1311 => data_o <= x"F4000029";
      when 1312 => data_o <= x"540002B4";
      when 1313 => data_o <= x"F4000DE3";
      when 1314 => data_o <= x"D2E7402B";
      when 1315 => data_o <= x"F4000DE3";
      when 1316 => data_o <= x"D27EC220";
      when 1317 => data_o <= x"F4000DDF";
      when 1318 => data_o <= x"D2E7402B";
      when 1319 => data_o <= x"F4000DDF";
      when 1320 => data_o <= x"D27EC220";
      when 1321 => data_o <= x"7400025D";
      when 1322 => data_o <= x"B9D0002B";
      when 1323 => data_o <= x"7400025D";
      when 1324 => data_o <= x"9FB08800";
      when 1325 => data_o <= x"F4000D0B";
      when 1326 => data_o <= x"D3D00040";
      when 1327 => data_o <= x"F4000000";
      when 1328 => data_o <= x"D1D0008D";
      when 1329 => data_o <= x"F4000D07";
      when 1330 => data_o <= x"D279C800";
      when 1331 => data_o <= x"F4000DD3";
      when 1332 => data_o <= x"D2EBBC9C";
      when 1333 => data_o <= x"7DD003ED";
      when 1334 => data_o <= x"04A3FC20";
      when 1335 => data_o <= x"74000077";
      when 1336 => data_o <= x"F4000D9D";
      when 1337 => data_o <= x"D36F4D08";
      when 1338 => data_o <= x"D0FEC800";
      when 1339 => data_o <= x"F4000D9F";
      when 1340 => data_o <= x"D0E7F628";
      when 1341 => data_o <= x"F4000D04";
      when 1342 => data_o <= x"D0FEC800";
      when 1343 => data_o <= x"F4000D00";
      when 1344 => data_o <= x"D0FEC220";
      when 1345 => data_o <= x"F4000D0B";
      when 1346 => data_o <= x"D01F4010";
      when 1347 => data_o <= x"0F6F401F";
      when 1348 => data_o <= x"4C97402B";
      when 1349 => data_o <= x"F4000010";
      when 1350 => data_o <= x"0DFF4DE3";
      when 1351 => data_o <= x"D2E48800";
      when 1352 => data_o <= x"7400024D";
      when 1353 => data_o <= x"F4000DE3";
      when 1354 => data_o <= x"D2EF400C";
      when 1355 => data_o <= x"0FD00DD3";
      when 1356 => data_o <= x"D2E9FB28";
      when 1357 => data_o <= x"F4000DE3";
      when 1358 => data_o <= x"D1500009";
      when 1359 => data_o <= x"F4000CFB";
      when 1360 => data_o <= x"D150000B";
      when 1361 => data_o <= x"F40012B8";
      when 1362 => data_o <= x"F40012BC";
      when 1363 => data_o <= x"7400052D";
      when 1364 => data_o <= x"7400026A";
      when 1365 => data_o <= x"54000541";
      when 1366 => data_o <= x"F4000DD3";
      when 1367 => data_o <= x"D2EB8308";
      when 1368 => data_o <= x"74000556";
      when 1369 => data_o <= x"5400023C";
      when 1370 => data_o <= x"D3D00007";
      when 1371 => data_o <= x"D1500558";
      when 1372 => data_o <= x"D3D00004";
      when 1373 => data_o <= x"54000558";
      when 1374 => data_o <= x"F4000004";
      when 1375 => data_o <= x"5400055A";
      when 1376 => data_o <= x"F4000008";
      when 1377 => data_o <= x"5400055A";
      when 1378 => data_o <= x"F4000080";
      when 1379 => data_o <= x"5400055C";
      when 1380 => data_o <= x"F4000001";
      when 1381 => data_o <= x"F4000DD7";
      when 1382 => data_o <= x"D27EC220";
      when 1383 => data_o <= x"F4000000";
      when 1384 => data_o <= x"F4000DD7";
      when 1385 => data_o <= x"D27EC220";
      when 1386 => data_o <= x"74000312";
      when 1387 => data_o <= x"740002A6";
      when 1388 => data_o <= x"F4000004";
      when 1389 => data_o <= x"74000556";
      when 1390 => data_o <= x"DBD00020";
      when 1391 => data_o <= x"4FA54572";
      when 1392 => data_o <= x"F4000020";
      when 1393 => data_o <= x"7400055C";
      when 1394 => data_o <= x"F4000DB3";
      when 1395 => data_o <= x"D3620000";
      when 1396 => data_o <= x"E9500580";
      when 1397 => data_o <= x"F4000000";
      when 1398 => data_o <= x"F4000DB3";
      when 1399 => data_o <= x"D0FEC800";
      when 1400 => data_o <= x"F4000DDF";
      when 1401 => data_o <= x"D2EF4003";
      when 1402 => data_o <= x"D1D00556";
      when 1403 => data_o <= x"7400004B";
      when 1404 => data_o <= x"D090D450";
      when 1405 => data_o <= x"D3D0FFFF";
      when 1406 => data_o <= x"4F4F400B";
      when 1407 => data_o <= x"D1D00558";
      when 1408 => data_o <= x"F4000000";
      when 1409 => data_o <= x"F4000DD7";
      when 1410 => data_o <= x"D27EC220";
      when 1411 => data_o <= x"7DD00525";
      when 1412 => data_o <= x"F4000DDF";
      when 1413 => data_o <= x"D2E28800";
      when 1414 => data_o <= x"7400052D";
      when 1415 => data_o <= x"F40000E0";
      when 1416 => data_o <= x"7400054F";
      when 1417 => data_o <= x"74000541";
      when 1418 => data_o <= x"F4000001";
      when 1419 => data_o <= x"F4000DB3";
      when 1420 => data_o <= x"D0FEC800";
      when 1421 => data_o <= x"54000564";
      when 1422 => data_o <= x"F40012AC";
      when 1423 => data_o <= x"54000583";
      when 1424 => data_o <= x"74000525";
      when 1425 => data_o <= x"740002A6";
      when 1426 => data_o <= x"F4000DDF";
      when 1427 => data_o <= x"D2E54564";
      when 1428 => data_o <= x"7400025D";
      when 1429 => data_o <= x"B8220000";
      when 1430 => data_o <= x"7400025D";
      when 1431 => data_o <= x"54000009";
      when 1432 => data_o <= x"7400025D";
      when 1433 => data_o <= x"BBC04800";
      when 1434 => data_o <= x"74000596";
      when 1435 => data_o <= x"54000093";
      when 1436 => data_o <= x"7400025D";
      when 1437 => data_o <= x"B9D00551";
      when 1438 => data_o <= x"54000596";
      when 1439 => data_o <= x"54000551";
      when 1440 => data_o <= x"74000529";
      when 1441 => data_o <= x"7400025D";
      when 1442 => data_o <= x"B9D00551";
      when 1443 => data_o <= x"F4000004";
      when 1444 => data_o <= x"54000598";
      when 1445 => data_o <= x"F4000DC7";
      when 1446 => data_o <= x"D2EF4DBF";
      when 1447 => data_o <= x"D27EC220";
      when 1448 => data_o <= x"54000302";
      when 1449 => data_o <= x"740003F7";
      when 1450 => data_o <= x"54000302";
      when 1451 => data_o <= x"54000312";
      when 1452 => data_o <= x"08800000";
      when 1453 => data_o <= x"F4000029";
      when 1454 => data_o <= x"740003DC";
      when 1455 => data_o <= x"EFB08800";
      when 1456 => data_o <= x"74000430";
      when 1457 => data_o <= x"54000302";
      when 1458 => data_o <= x"F4000008";
      when 1459 => data_o <= x"D090C184";
      when 1460 => data_o <= x"7400004B";
      when 1461 => data_o <= x"F150004B";
      when 1462 => data_o <= x"740005B2";
      when 1463 => data_o <= x"F40012A4";
      when 1464 => data_o <= x"6E4D0426";
      when 1465 => data_o <= x"7400040B";
      when 1466 => data_o <= x"07A545BC";
      when 1467 => data_o <= x"540005B6";
      when 1468 => data_o <= x"EFB08800";
      when 1469 => data_o <= x"7400042C";
      when 1470 => data_o <= x"740005B2";
      when 1471 => data_o <= x"F40012A4";
      when 1472 => data_o <= x"6E420000";
      when 1473 => data_o <= x"E95005C3";
      when 1474 => data_o <= x"5400030B";
      when 1475 => data_o <= x"74000302";
      when 1476 => data_o <= x"F4000C2C";
      when 1477 => data_o <= x"5400030B";
      when 1478 => data_o <= x"F4000003";
      when 1479 => data_o <= x"D1D00556";
      when 1480 => data_o <= x"7400004B";
      when 1481 => data_o <= x"5400030B";
      when 1482 => data_o <= x"F4000DD7";
      when 1483 => data_o <= x"D2E93D0D";
      when 1484 => data_o <= x"D135410E";
      when 1485 => data_o <= x"740005CA";
      when 1486 => data_o <= x"F4000DDF";
      when 1487 => data_o <= x"D2EF0800";
      when 1488 => data_o <= x"F400FA00";
      when 1489 => data_o <= x"74000070";
      when 1490 => data_o <= x"E95005D4";
      when 1491 => data_o <= x"84924800";
      when 1492 => data_o <= x"F4000DB5";
      when 1493 => data_o <= x"D3674070";
      when 1494 => data_o <= x"E95005D8";
      when 1495 => data_o <= x"740002A6";
      when 1496 => data_o <= x"F4000DDF";
      when 1497 => data_o <= x"D2E08800";
      when 1498 => data_o <= x"F4000015";
      when 1499 => data_o <= x"540002C5";
      when 1500 => data_o <= x"F4000DB5";
      when 1501 => data_o <= x"D36F4000";
      when 1502 => data_o <= x"D397409D";
      when 1503 => data_o <= x"D1D005DA";
      when 1504 => data_o <= x"F4000018";
      when 1505 => data_o <= x"7400009D";
      when 1506 => data_o <= x"0FD00060";
      when 1507 => data_o <= x"94000000";
      when 1508 => data_o <= x"0C220000";
      when 1509 => data_o <= x"740005CA";
      when 1510 => data_o <= x"740002A6";
      when 1511 => data_o <= x"04800000";
      when 1512 => data_o <= x"F4FFFFFF";
      when 1513 => data_o <= x"4FCF4018";
      when 1514 => data_o <= x"740000A2";
      when 1515 => data_o <= x"07D0001F";
      when 1516 => data_o <= x"4FCF4005";
      when 1517 => data_o <= x"740000A2";
      when 1518 => data_o <= x"F4000003";
      when 1519 => data_o <= x"6E493D15";
      when 1520 => data_o <= x"D137410E";
      when 1521 => data_o <= x"F4000000";
      when 1522 => data_o <= x"D3C7409D";
      when 1523 => data_o <= x"F4000DDF";
      when 1524 => data_o <= x"D2E71C0C";
      when 1525 => data_o <= x"F150023C";
      when 1526 => data_o <= x"740005CA";
      when 1527 => data_o <= x"740002A6";
      when 1528 => data_o <= x"F4000DDF";
      when 1529 => data_o <= x"D2EF4040";
      when 1530 => data_o <= x"94000000";
      when 1531 => data_o <= x"0C220000";
      when 1532 => data_o <= x"740005CA";
      when 1533 => data_o <= x"51407D38";
      when 1534 => data_o <= x"94000000";
      when 1535 => data_o <= x"4FD00010";
      when 1536 => data_o <= x"94000000";
      when 1537 => data_o <= x"6E493D15";
      when 1538 => data_o <= x"D137410E";
      when 1539 => data_o <= x"F43FFFFF";
      when 1540 => data_o <= x"4D5005DA";
      when 1541 => data_o <= x"F400000E";
      when 1542 => data_o <= x"740005CD";
      when 1543 => data_o <= x"540005DC";
      when 1544 => data_o <= x"F4000014";
      when 1545 => data_o <= x"740005CD";
      when 1546 => data_o <= x"F4000038";
      when 1547 => data_o <= x"740002B4";
      when 1548 => data_o <= x"540005DC";
      when 1549 => data_o <= x"F4000014";
      when 1550 => data_o <= x"740005CD";
      when 1551 => data_o <= x"F400003A";
      when 1552 => data_o <= x"740002B4";
      when 1553 => data_o <= x"540005DC";
      when 1554 => data_o <= x"F4000014";
      when 1555 => data_o <= x"740005CD";
      when 1556 => data_o <= x"F4000030";
      when 1557 => data_o <= x"740002B4";
      when 1558 => data_o <= x"540005DC";
      when 1559 => data_o <= x"74000605";
      when 1560 => data_o <= x"F15005E5";
      when 1561 => data_o <= x"740005CA";
      when 1562 => data_o <= x"7DD0060D";
      when 1563 => data_o <= x"28220000";
      when 1564 => data_o <= x"740005CA";
      when 1565 => data_o <= x"7DD00612";
      when 1566 => data_o <= x"28220000";
      when 1567 => data_o <= x"740005FC";
      when 1568 => data_o <= x"540005E5";
      when 1569 => data_o <= x"F4000014";
      when 1570 => data_o <= x"740005CD";
      when 1571 => data_o <= x"EFD00030";
      when 1572 => data_o <= x"740002B4";
      when 1573 => data_o <= x"540005FC";
      when 1574 => data_o <= x"F4000014";
      when 1575 => data_o <= x"740005CD";
      when 1576 => data_o <= x"EFD0003A";
      when 1577 => data_o <= x"740002B4";
      when 1578 => data_o <= x"540005FC";
      when 1579 => data_o <= x"740005F6";
      when 1580 => data_o <= x"F4000190";
      when 1581 => data_o <= x"7400030B";
      when 1582 => data_o <= x"54000605";
      when 1583 => data_o <= x"F400001F";
      when 1584 => data_o <= x"740002B4";
      when 1585 => data_o <= x"5400062B";
      when 1586 => data_o <= x"F1D005FC";
      when 1587 => data_o <= x"540005E5";
      when 1588 => data_o <= x"F4000DDF";
      when 1589 => data_o <= x"D2EF52AC";
      when 1590 => data_o <= x"7400052D";
      when 1591 => data_o <= x"07D00D0B";
      when 1592 => data_o <= x"D173FB20";
      when 1593 => data_o <= x"F40000C0";
      when 1594 => data_o <= x"7400054F";
      when 1595 => data_o <= x"74000541";
      when 1596 => data_o <= x"540002A6";
      when 1597 => data_o <= x"F4000001";
      when 1598 => data_o <= x"74000634";
      when 1599 => data_o <= x"F4000003";
      when 1600 => data_o <= x"94FFFFFF";
      when 1601 => data_o <= x"F4000015";
      when 1602 => data_o <= x"540002C5";
      when 1603 => data_o <= x"514F4004";
      when 1604 => data_o <= x"94000000";
      when 1605 => data_o <= x"D090C800";
      when 1606 => data_o <= x"74000430";
      when 1607 => data_o <= x"5400023C";
      when 1608 => data_o <= x"F4000002";
      when 1609 => data_o <= x"74000634";
      when 1610 => data_o <= x"74000529";
      when 1611 => data_o <= x"74000594";
      when 1612 => data_o <= x"F4000D9C";
      when 1613 => data_o <= x"D36F4001";
      when 1614 => data_o <= x"6E4F4008";
      when 1615 => data_o <= x"4C374302";
      when 1616 => data_o <= x"F4000002";
      when 1617 => data_o <= x"740002B4";
      when 1618 => data_o <= x"F4000DA7";
      when 1619 => data_o <= x"D2EF403F";
      when 1620 => data_o <= x"D3D00DB5";
      when 1621 => data_o <= x"D367409D";
      when 1622 => data_o <= x"D0374268";
      when 1623 => data_o <= x"540002A7";
      when 1624 => data_o <= x"BBD000FC";
      when 1625 => data_o <= x"94000000";
      when 1626 => data_o <= x"4FD000D0";
      when 1627 => data_o <= x"94000000";
      when 1628 => data_o <= x"6E408800";
      when 1629 => data_o <= x"9BDFFFFF";
      when 1630 => data_o <= x"4FC06E7C";
      when 1631 => data_o <= x"74000658";
      when 1632 => data_o <= x"E9500663";
      when 1633 => data_o <= x"D0AF7FFF";
      when 1634 => data_o <= x"54000664";
      when 1635 => data_o <= x"2BDFFFFF";
      when 1636 => data_o <= x"05F4C128";
      when 1637 => data_o <= x"6E408800";
      when 1638 => data_o <= x"7400065D";
      when 1639 => data_o <= x"EFB08800";
      when 1640 => data_o <= x"29453D03";
      when 1641 => data_o <= x"D1D00556";
      when 1642 => data_o <= x"7400004B";
      when 1643 => data_o <= x"8417C800";
      when 1644 => data_o <= x"74000658";
      when 1645 => data_o <= x"E9500671";
      when 1646 => data_o <= x"F42ABFFF";
      when 1647 => data_o <= x"D0800000";
      when 1648 => data_o <= x"54000673";
      when 1649 => data_o <= x"F40000F5";
      when 1650 => data_o <= x"94500000";
      when 1651 => data_o <= x"0CA5423C";
      when 1652 => data_o <= x"F4000000";
      when 1653 => data_o <= x"08800000";
      when 1654 => data_o <= x"F4000184";
      when 1655 => data_o <= x"7400030B";
      when 1656 => data_o <= x"54000605";
      when 1657 => data_o <= x"54000617";
      when 1658 => data_o <= x"F4001378";
      when 1659 => data_o <= x"7400030B";
      when 1660 => data_o <= x"74000022";
      when 1661 => data_o <= x"E9500680";
      when 1662 => data_o <= x"740005E5";
      when 1663 => data_o <= x"5400067C";
      when 1664 => data_o <= x"08800000";
      when 1665 => data_o <= x"740005CA";
      when 1666 => data_o <= x"740002A6";
      when 1667 => data_o <= x"F400003C";
      when 1668 => data_o <= x"740002B4";
      when 1669 => data_o <= x"F4000034";
      when 1670 => data_o <= x"740002B4";
      when 1671 => data_o <= x"F4000009";
      when 1672 => data_o <= x"740002B4";
      when 1673 => data_o <= x"F400001F";
      when 1674 => data_o <= x"740002B4";
      when 1675 => data_o <= x"F400001F";
      when 1676 => data_o <= x"740002B4";
      when 1677 => data_o <= x"740005F6";
      when 1678 => data_o <= x"F4000000";
      when 1679 => data_o <= x"F4000D0B";
      when 1680 => data_o <= x"D27EC220";
      when 1681 => data_o <= x"740005CA";
      when 1682 => data_o <= x"F4000138";
      when 1683 => data_o <= x"7400030B";
      when 1684 => data_o <= x"74000605";
      when 1685 => data_o <= x"F4000004";
      when 1686 => data_o <= x"F4000D0B";
      when 1687 => data_o <= x"D279FB20";
      when 1688 => data_o <= x"540005F6";
      when 1689 => data_o <= x"F4000D0B";
      when 1690 => data_o <= x"D017E604";
      when 1691 => data_o <= x"84A9FB0C";
      when 1692 => data_o <= x"9FB08800";
      when 1693 => data_o <= x"F4000D0B";
      when 1694 => data_o <= x"D0106E0C";
      when 1695 => data_o <= x"B9FF4003";
      when 1696 => data_o <= x"D3C74009";
      when 1697 => data_o <= x"28220000";
      when 1698 => data_o <= x"740005CA";
      when 1699 => data_o <= x"F400017C";
      when 1700 => data_o <= x"7400030B";
      when 1701 => data_o <= x"74000605";
      when 1702 => data_o <= x"54000699";
      when 1703 => data_o <= x"F4000D0B";
      when 1704 => data_o <= x"D2E20000";
      when 1705 => data_o <= x"E95006AD";
      when 1706 => data_o <= x"7400069D";
      when 1707 => data_o <= x"740005E5";
      when 1708 => data_o <= x"540006A7";
      when 1709 => data_o <= x"08800000";
      when 1710 => data_o <= x"740005CA";
      when 1711 => data_o <= x"F400014C";
      when 1712 => data_o <= x"7400030B";
      when 1713 => data_o <= x"740005FC";
      when 1714 => data_o <= x"540006A7";
      when 1715 => data_o <= x"740005CA";
      when 1716 => data_o <= x"F400015C";
      when 1717 => data_o <= x"7400030B";
      when 1718 => data_o <= x"740005FC";
      when 1719 => data_o <= x"540006A7";
      when 1720 => data_o <= x"740005CA";
      when 1721 => data_o <= x"F4000012";
      when 1722 => data_o <= x"540002B4";
      when 1723 => data_o <= x"F4000022";
      when 1724 => data_o <= x"740003DC";
      when 1725 => data_o <= x"05F74279";
      when 1726 => data_o <= x"F4000DDF";
      when 1727 => data_o <= x"D2E48800";
      when 1728 => data_o <= x"7400024D";
      when 1729 => data_o <= x"2BD00DDF";
      when 1730 => data_o <= x"D1500009";
      when 1731 => data_o <= x"F400019C";
      when 1732 => data_o <= x"7400030B";
      when 1733 => data_o <= x"740006BB";
      when 1734 => data_o <= x"54000525";
      when 1735 => data_o <= x"740006C3";
      when 1736 => data_o <= x"F400000E";
      when 1737 => data_o <= x"740002B4";
      when 1738 => data_o <= x"F40004B0";
      when 1739 => data_o <= x"5400030B";
      when 1740 => data_o <= x"F4000000";
      when 1741 => data_o <= x"D150010E";
      when 1742 => data_o <= x"7400060D";
      when 1743 => data_o <= x"740006C7";
      when 1744 => data_o <= x"F4001B30";
      when 1745 => data_o <= x"7400030B";
      when 1746 => data_o <= x"540005E5";
      when 1747 => data_o <= x"F4000022";
      when 1748 => data_o <= x"740003DC";
      when 1749 => data_o <= x"F4000DDB";
      when 1750 => data_o <= x"D2EF4080";
      when 1751 => data_o <= x"0C17F9F0";
      when 1752 => data_o <= x"3FC74077";
      when 1753 => data_o <= x"28220000";
      when 1754 => data_o <= x"740006C3";
      when 1755 => data_o <= x"F400000E";
      when 1756 => data_o <= x"540002B4";
      when 1757 => data_o <= x"740006D3";
      when 1758 => data_o <= x"38220000";
      when 1759 => data_o <= x"540006D3";
      when 1760 => data_o <= x"F4000DC7";
      when 1761 => data_o <= x"D150002D";
      when 1762 => data_o <= x"F4000DCB";
      when 1763 => data_o <= x"D3D00005";
      when 1764 => data_o <= x"05F7C800";
      when 1765 => data_o <= x"74000064";
      when 1766 => data_o <= x"540006E8";
      when 1767 => data_o <= x"9BC546E5";
      when 1768 => data_o <= x"ECA08800";
      when 1769 => data_o <= x"F4000005";
      when 1770 => data_o <= x"E5B92420";
      when 1771 => data_o <= x"F400003E";
      when 1772 => data_o <= x"D137410E";
      when 1773 => data_o <= x"F4000DCB";
      when 1774 => data_o <= x"D391040C";
      when 1775 => data_o <= x"F1F20000";
      when 1776 => data_o <= x"74000064";
      when 1777 => data_o <= x"540006F5";
      when 1778 => data_o <= x"F4000004";
      when 1779 => data_o <= x"D090FCE4";
      when 1780 => data_o <= x"9FB546F0";
      when 1781 => data_o <= x"05B08800";
      when 1782 => data_o <= x"740006E2";
      when 1783 => data_o <= x"7400039B";
      when 1784 => data_o <= x"F4000DC7";
      when 1785 => data_o <= x"D279FBF4";
      when 1786 => data_o <= x"F4000DBF";
      when 1787 => data_o <= x"D27EFD00";
      when 1788 => data_o <= x"D3D00DCB";
      when 1789 => data_o <= x"D27EC800";
      when 1790 => data_o <= x"F400121C";
      when 1791 => data_o <= x"74000106";
      when 1792 => data_o <= x"04800000";
      when 1793 => data_o <= x"E9500707";
      when 1794 => data_o <= x"74000148";
      when 1795 => data_o <= x"740006E0";
      when 1796 => data_o <= x"7400012C";
      when 1797 => data_o <= x"74000148";
      when 1798 => data_o <= x"74000567";
      when 1799 => data_o <= x"740003A1";
      when 1800 => data_o <= x"740006E9";
      when 1801 => data_o <= x"ED50010E";
      when 1802 => data_o <= x"7400003F";
      when 1803 => data_o <= x"74000022";
      when 1804 => data_o <= x"E9500711";
      when 1805 => data_o <= x"F4000000";
      when 1806 => data_o <= x"7400018B";
      when 1807 => data_o <= x"F400007C";
      when 1808 => data_o <= x"74000146";
      when 1809 => data_o <= x"74000067";
      when 1810 => data_o <= x"3E6B6F03";
      when 1811 => data_o <= x"39D0012C";
      when 1812 => data_o <= x"F4000D93";
      when 1813 => data_o <= x"D3D00088";
      when 1814 => data_o <= x"740001A8";
      when 1815 => data_o <= x"F4000DC7";
      when 1816 => data_o <= x"D27EFD00";
      when 1817 => data_o <= x"F4000DBF";
      when 1818 => data_o <= x"D27EC800";
      when 1819 => data_o <= x"74000148";
      when 1820 => data_o <= x"F4000000";
      when 1821 => data_o <= x"08800000";
      when 1822 => data_o <= x"7400070A";
      when 1823 => data_o <= x"EDD00487";
      when 1824 => data_o <= x"5400071E";
      when 1825 => data_o <= x"08800000";
      when 1826 => data_o <= x"74000148";
      when 1827 => data_o <= x"74000067";
      when 1828 => data_o <= x"72724506";
      when 1829 => data_o <= x"FF23726F";
      when 1830 => data_o <= x"39D0012C";
      when 1831 => data_o <= x"74000192";
      when 1832 => data_o <= x"74000148";
      when 1833 => data_o <= x"F4000D93";
      when 1834 => data_o <= x"D3D00DC7";
      when 1835 => data_o <= x"D2E7412C";
      when 1836 => data_o <= x"54000148";
      when 1837 => data_o <= x"F4000000";
      when 1838 => data_o <= x"A7FF4008";
      when 1839 => data_o <= x"A6EF4004";
      when 1840 => data_o <= x"D090EF20";
      when 1841 => data_o <= x"F4000D93";
      when 1842 => data_o <= x"D3D00DC3";
      when 1843 => data_o <= x"D27EFD00";
      when 1844 => data_o <= x"07D00DD7";
      when 1845 => data_o <= x"D27EC120";
      when 1846 => data_o <= x"F4000DB3";
      when 1847 => data_o <= x"D27EC800";
      when 1848 => data_o <= x"F4000DBB";
      when 1849 => data_o <= x"D27EC800";
      when 1850 => data_o <= x"F4001C78";
      when 1851 => data_o <= x"74000106";
      when 1852 => data_o <= x"74000022";
      when 1853 => data_o <= x"E950073F";
      when 1854 => data_o <= x"74000722";
      when 1855 => data_o <= x"F400000C";
      when 1856 => data_o <= x"A6EDC800";
      when 1857 => data_o <= x"5400072D";
      when 1858 => data_o <= x"08800000";
      when 1859 => data_o <= x"F4000DDB";
      when 1860 => data_o <= x"D017EE04";
      when 1861 => data_o <= x"84A9FB7C";
      when 1862 => data_o <= x"F4000000";
      when 1863 => data_o <= x"4A7EFD12";
      when 1864 => data_o <= x"94345678";
      when 1865 => data_o <= x"7400026A";
      when 1866 => data_o <= x"04800000";
      when 1867 => data_o <= x"E9500757";
      when 1868 => data_o <= x"48800000";
      when 1869 => data_o <= x"F5000000";
      when 1870 => data_o <= x"D090C800";
      when 1871 => data_o <= x"7400026A";
      when 1872 => data_o <= x"05D0027B";
      when 1873 => data_o <= x"D0920000";
      when 1874 => data_o <= x"7CE7427B";
      when 1875 => data_o <= x"28920000";
      when 1876 => data_o <= x"C1500752";
      when 1877 => data_o <= x"EFB28800";
      when 1878 => data_o <= x"54000521";
      when 1879 => data_o <= x"EFB28120";
      when 1880 => data_o <= x"5400026A";
      when 1881 => data_o <= x"F4000000";
      when 1882 => data_o <= x"05500743";
      when 1883 => data_o <= x"06C20000";
      when 1884 => data_o <= x"E9500761";
      when 1885 => data_o <= x"ECEF401F";
      when 1886 => data_o <= x"4DD0012C";
      when 1887 => data_o <= x"74000156";
      when 1888 => data_o <= x"54000764";
      when 1889 => data_o <= x"F4000003";
      when 1890 => data_o <= x"740001A0";
      when 1891 => data_o <= x"EC800000";
      when 1892 => data_o <= x"08800000";
      when 1893 => data_o <= x"04800000";
      when 1894 => data_o <= x"F1D0004B";
      when 1895 => data_o <= x"06420000";
      when 1896 => data_o <= x"E9500766";
      when 1897 => data_o <= x"EFD00010";
      when 1898 => data_o <= x"D090C800";
      when 1899 => data_o <= x"06EF4012";
      when 1900 => data_o <= x"94345678";
      when 1901 => data_o <= x"6E490800";
      when 1902 => data_o <= x"E9500771";
      when 1903 => data_o <= x"D21D0800";
      when 1904 => data_o <= x"5400076B";
      when 1905 => data_o <= x"8665475B";
      when 1906 => data_o <= x"04E74419";
      when 1907 => data_o <= x"E4800000";
      when 1908 => data_o <= x"E9500776";
      when 1909 => data_o <= x"EC16C220";
      when 1910 => data_o <= x"7FBECA20";
      when 1911 => data_o <= x"540005B6";
      when 1912 => data_o <= x"F4000DB7";
      when 1913 => data_o <= x"D367C800";
      when 1914 => data_o <= x"74000064";
      when 1915 => data_o <= x"54000780";
      when 1916 => data_o <= x"48410800";
      when 1917 => data_o <= x"F4000D9B";
      when 1918 => data_o <= x"D03B8800";
      when 1919 => data_o <= x"5400077A";
      when 1920 => data_o <= x"F4000DB7";
      when 1921 => data_o <= x"D3608800";
      when 1922 => data_o <= x"06C20000";
      when 1923 => data_o <= x"E9500786";
      when 1924 => data_o <= x"EFD00CCB";
      when 1925 => data_o <= x"D3D00001";
      when 1926 => data_o <= x"07D00DB7";
      when 1927 => data_o <= x"D0FEFD00";
      when 1928 => data_o <= x"7400004E";
      when 1929 => data_o <= x"5400078F";
      when 1930 => data_o <= x"48410800";
      when 1931 => data_o <= x"F4000D9B";
      when 1932 => data_o <= x"D039FB20";
      when 1933 => data_o <= x"74000053";
      when 1934 => data_o <= x"5400078A";
      when 1935 => data_o <= x"08800000";
      when 1936 => data_o <= x"F4000DD3";
      when 1937 => data_o <= x"D27EC220";
      when 1938 => data_o <= x"F4000DD3";
      when 1939 => data_o <= x"D2E08800";
      when 1940 => data_o <= x"F4000000";
      when 1941 => data_o <= x"D1500782";
      when 1942 => data_o <= x"74000778";
      when 1943 => data_o <= x"E7C24800";
      when 1944 => data_o <= x"54000782";
      when 1945 => data_o <= x"74000778";
      when 1946 => data_o <= x"F3BD09D0";
      when 1947 => data_o <= x"54000782";
      when 1948 => data_o <= x"74000778";
      when 1949 => data_o <= x"E5D00790";
      when 1950 => data_o <= x"54000782";
      when 1951 => data_o <= x"F4000CCB";
      when 1952 => data_o <= x"D01F4001";
      when 1953 => data_o <= x"74000782";
      when 1954 => data_o <= x"54000790";
      when 1955 => data_o <= x"74000778";
      when 1956 => data_o <= x"F3BF4CCB";
      when 1957 => data_o <= x"D3C54782";
      when 1958 => data_o <= x"74000067";
      when 1959 => data_o <= x"6F43200A";
      when 1960 => data_o <= x"7865746E";
      when 1961 => data_o <= x"FF203A74";
      when 1962 => data_o <= x"39D0012C";
      when 1963 => data_o <= x"F4000D9B";
      when 1964 => data_o <= x"D3D00DB7";
      when 1965 => data_o <= x"D36F4000";
      when 1966 => data_o <= x"7400004E";
      when 1967 => data_o <= x"540007B3";
      when 1968 => data_o <= x"99D00765";
      when 1969 => data_o <= x"74000053";
      when 1970 => data_o <= x"540007B0";
      when 1971 => data_o <= x"EDD00148";
      when 1972 => data_o <= x"74000067";
      when 1973 => data_o <= x"7543200A";
      when 1974 => data_o <= x"6E657272";
      when 1975 => data_o <= x"FF203A74";
      when 1976 => data_o <= x"39D0012C";
      when 1977 => data_o <= x"F4000DD3";
      when 1978 => data_o <= x"D2E74765";
      when 1979 => data_o <= x"54000148";
      when 1980 => data_o <= x"04800000";
      when 1981 => data_o <= x"EBBEFB08";
      when 1982 => data_o <= x"7400003B";
      when 1983 => data_o <= x"E95007C8";
      when 1984 => data_o <= x"7400003D";
      when 1985 => data_o <= x"E5D0001F";
      when 1986 => data_o <= x"740003F9";
      when 1987 => data_o <= x"E95007C5";
      when 1988 => data_o <= x"EFBEC220";
      when 1989 => data_o <= x"EFB7DFF5";
      when 1990 => data_o <= x"740000E6";
      when 1991 => data_o <= x"28A547BE";
      when 1992 => data_o <= x"EFBEC16E";
      when 1993 => data_o <= x"B8800000";
      when 1994 => data_o <= x"05F84E04";
      when 1995 => data_o <= x"7FD0001F";
      when 1996 => data_o <= x"4DD0001F";
      when 1997 => data_o <= x"7400001F";
      when 1998 => data_o <= x"7400001D";
      when 1999 => data_o <= x"740007BC";
      when 2000 => data_o <= x"E95007DF";
      when 2001 => data_o <= x"292F4008";
      when 2002 => data_o <= x"D090DD4B";
      when 2003 => data_o <= x"F40012A4";
      when 2004 => data_o <= x"6E420000";
      when 2005 => data_o <= x"E95007D8";
      when 2006 => data_o <= x"F4000020";
      when 2007 => data_o <= x"0C800000";
      when 2008 => data_o <= x"F4000005";
      when 2009 => data_o <= x"740000A2";
      when 2010 => data_o <= x"7400035B";
      when 2011 => data_o <= x"7400012C";
      when 2012 => data_o <= x"7400033E";
      when 2013 => data_o <= x"74000156";
      when 2014 => data_o <= x"540007E0";
      when 2015 => data_o <= x"2BBEFB20";
      when 2016 => data_o <= x"29D0004B";
      when 2017 => data_o <= x"06420000";
      when 2018 => data_o <= x"E95007CA";
      when 2019 => data_o <= x"ED500148";
      when 2020 => data_o <= x"740003ED";
      when 2021 => data_o <= x"F4000DB7";
      when 2022 => data_o <= x"D3620000";
      when 2023 => data_o <= x"D09D0800";
      when 2024 => data_o <= x"C15007EE";
      when 2025 => data_o <= x"05F10420";
      when 2026 => data_o <= x"F4000D9B";
      when 2027 => data_o <= x"D03B8800";
      when 2028 => data_o <= x"740007C9";
      when 2029 => data_o <= x"295007E7";
      when 2030 => data_o <= x"EFBEC220";
      when 2031 => data_o <= x"740003ED";
      when 2032 => data_o <= x"540007C9";
      when 2033 => data_o <= x"64032E01";
      when 2034 => data_o <= x"65047075";
      when 2035 => data_o <= x"01746978";
      when 2036 => data_o <= x"2A32022B";
      when 2037 => data_o <= x"3F013F01";
      when 2038 => data_o <= x"5F013F01";
      when 2039 => data_o <= x"022B3102";
      when 2040 => data_o <= x"3F013E72";
      when 2041 => data_o <= x"632A3203";
      when 2042 => data_o <= x"65737504";
      when 2043 => data_o <= x"40630372";
      when 2044 => data_o <= x"2163032B";
      when 2045 => data_o <= x"023F012B";
      when 2046 => data_o <= x"72027072";
      when 2047 => data_o <= x"6E610340";
      when 2048 => data_o <= x"2F320264";
      when 2049 => data_o <= x"706D6A03";
      when 2050 => data_o <= x"2B407703";
      when 2051 => data_o <= x"2B217703";
      when 2052 => data_o <= x"73023F01";
      when 2053 => data_o <= x"033F0170";
      when 2054 => data_o <= x"03726F78";
      when 2055 => data_o <= x"042F3275";
      when 2056 => data_o <= x"6C6C6163";
      when 2057 => data_o <= x"02407702";
      when 2058 => data_o <= x"7205723E";
      when 2059 => data_o <= x"63747065";
      when 2060 => data_o <= x"012B3402";
      when 2061 => data_o <= x"2B63023F";
      when 2062 => data_o <= x"043D3002";
      when 2063 => data_o <= x"7874696C";
      when 2064 => data_o <= x"022B4002";
      when 2065 => data_o <= x"2D052B21";
      when 2066 => data_o <= x"74706572";
      when 2067 => data_o <= x"01707502";
      when 2068 => data_o <= x"023F013F";
      when 2069 => data_o <= x"40033C30";
      when 2070 => data_o <= x"40017361";
      when 2071 => data_o <= x"21707203";
      when 2072 => data_o <= x"66692D04";
      when 2073 => data_o <= x"6F70043A";
      when 2074 => data_o <= x"3F017472";
      when 2075 => data_o <= x"63033F01";
      when 2076 => data_o <= x"21036D6F";
      when 2077 => data_o <= x"63027361";
      when 2078 => data_o <= x"70730340";
      when 2079 => data_o <= x"66690421";
      when 2080 => data_o <= x"6F043A63";
      when 2081 => data_o <= x"04726576";
      when 2082 => data_o <= x"3A7A6669";
      when 2083 => data_o <= x"6F726404";
      when 2084 => data_o <= x"77730470";
      when 2085 => data_o <= x"6C037061";
      when 2086 => data_o <= x"3F017469";
      when 2087 => data_o <= x"21707503";
      when 2088 => data_o <= x"F4001FC4";
      when 2089 => data_o <= x"E4800000";
      when 2090 => data_o <= x"E950082D";
      when 2091 => data_o <= x"383F3424";
      when 2092 => data_o <= x"D3C54829";
      when 2093 => data_o <= x"F3B38220";
      when 2094 => data_o <= x"0D151D07";
      when 2095 => data_o <= x"352D253D";
      when 2096 => data_o <= x"FF151D02";
      when 2097 => data_o <= x"F1F38800";
      when 2098 => data_o <= x"04800000";
      when 2099 => data_o <= x"E950083A";
      when 2100 => data_o <= x"F0E49B90";
      when 2101 => data_o <= x"E9500838";
      when 2102 => data_o <= x"2BBEFBF5";
      when 2103 => data_o <= x"08800000";
      when 2104 => data_o <= x"F3427420";
      when 2105 => data_o <= x"54000832";
      when 2106 => data_o <= x"2BBF3B08";
      when 2107 => data_o <= x"E7487420";
      when 2108 => data_o <= x"7400004B";
      when 2109 => data_o <= x"E5B90800";
      when 2110 => data_o <= x"E9500840";
      when 2111 => data_o <= x"EE104220";
      when 2112 => data_o <= x"F1D0004B";
      when 2113 => data_o <= x"F3990800";
      when 2114 => data_o <= x"E950083B";
      when 2115 => data_o <= x"F0220000";
      when 2116 => data_o <= x"F4000DB7";
      when 2117 => data_o <= x"D3620000";
      when 2118 => data_o <= x"04800000";
      when 2119 => data_o <= x"E9500851";
      when 2120 => data_o <= x"D09D017C";
      when 2121 => data_o <= x"104F4D9B";
      when 2122 => data_o <= x"D03B9D4B";
      when 2123 => data_o <= x"E5D0083B";
      when 2124 => data_o <= x"E9500850";
      when 2125 => data_o <= x"2BBF3B38";
      when 2126 => data_o <= x"F400001F";
      when 2127 => data_o <= x"4C220000";
      when 2128 => data_o <= x"ECA54846";
      when 2129 => data_o <= x"08800000";
      when 2130 => data_o <= x"05FF60B8";
      when 2131 => data_o <= x"74000831";
      when 2132 => data_o <= x"E9500869";
      when 2133 => data_o <= x"E79F4000";
      when 2134 => data_o <= x"D3C7409D";
      when 2135 => data_o <= x"D1348800";
      when 2136 => data_o <= x"F40020C0";
      when 2137 => data_o <= x"74000831";
      when 2138 => data_o <= x"E9500866";
      when 2139 => data_o <= x"10474844";
      when 2140 => data_o <= x"04800000";
      when 2141 => data_o <= x"E9500862";
      when 2142 => data_o <= x"7400034D";
      when 2143 => data_o <= x"7400012C";
      when 2144 => data_o <= x"74000156";
      when 2145 => data_o <= x"54000865";
      when 2146 => data_o <= x"EDD00353";
      when 2147 => data_o <= x"F4000003";
      when 2148 => data_o <= x"740001A0";
      when 2149 => data_o <= x"54000868";
      when 2150 => data_o <= x"74000350";
      when 2151 => data_o <= x"74000192";
      when 2152 => data_o <= x"EFD00005";
      when 2153 => data_o <= x"29D00828";
      when 2154 => data_o <= x"74000356";
      when 2155 => data_o <= x"7400012C";
      when 2156 => data_o <= x"74000156";
      when 2157 => data_o <= x"F4000006";
      when 2158 => data_o <= x"D090C220";
      when 2159 => data_o <= x"F400001A";
      when 2160 => data_o <= x"06C90800";
      when 2161 => data_o <= x"E9500876";
      when 2162 => data_o <= x"E79740A2";
      when 2163 => data_o <= x"F400003F";
      when 2164 => data_o <= x"4DD00852";
      when 2165 => data_o <= x"54000870";
      when 2166 => data_o <= x"E7D00003";
      when 2167 => data_o <= x"4F9F4003";
      when 2168 => data_o <= x"D1B90800";
      when 2169 => data_o <= x"E950087C";
      when 2170 => data_o <= x"74000852";
      when 2171 => data_o <= x"04800000";
      when 2172 => data_o <= x"EFBEC800";
      when 2173 => data_o <= x"5400033E";
      when 2174 => data_o <= x"05F74347";
      when 2175 => data_o <= x"07D00003";
      when 2176 => data_o <= x"740001A0";
      when 2177 => data_o <= x"99D00356";
      when 2178 => data_o <= x"07D00007";
      when 2179 => data_o <= x"740001A0";
      when 2180 => data_o <= x"7400086F";
      when 2181 => data_o <= x"29D00844";
      when 2182 => data_o <= x"04800000";
      when 2183 => data_o <= x"E950088E";
      when 2184 => data_o <= x"74000067";
      when 2185 => data_o <= x"FF205C02";
      when 2186 => data_o <= x"39D0012C";
      when 2187 => data_o <= x"7400034A";
      when 2188 => data_o <= x"7400012C";
      when 2189 => data_o <= x"5400088F";
      when 2190 => data_o <= x"EFB20000";
      when 2191 => data_o <= x"7400033E";
      when 2192 => data_o <= x"54000148";
      when 2193 => data_o <= x"E6E07D1A";
      when 2194 => data_o <= x"740000A2";
      when 2195 => data_o <= x"F4000015";
      when 2196 => data_o <= x"6E420000";
      when 2197 => data_o <= x"E9500899";
      when 2198 => data_o <= x"F3B20000";
      when 2199 => data_o <= x"F7FFFFFF";
      when 2200 => data_o <= x"4C410108";
      when 2201 => data_o <= x"05B08800";
      when 2202 => data_o <= x"07D00001";
      when 2203 => data_o <= x"6E420000";
      when 2204 => data_o <= x"E95008A9";
      when 2205 => data_o <= x"74000891";
      when 2206 => data_o <= x"E95008A9";
      when 2207 => data_o <= x"F1D0087E";
      when 2208 => data_o <= x"EFD0000A";
      when 2209 => data_o <= x"F400000E";
      when 2210 => data_o <= x"74000158";
      when 2211 => data_o <= x"74000067";
      when 2212 => data_o <= x"6665720A";
      when 2213 => data_o <= x"20737265";
      when 2214 => data_o <= x"FF3A6F74";
      when 2215 => data_o <= x"39D0012C";
      when 2216 => data_o <= x"74000148";
      when 2217 => data_o <= x"04800000";
      when 2218 => data_o <= x"E95008AE";
      when 2219 => data_o <= x"7DD0087E";
      when 2220 => data_o <= x"2B427420";
      when 2221 => data_o <= x"540008A9";
      when 2222 => data_o <= x"EFB08800";
      when 2223 => data_o <= x"7400042C";
      when 2224 => data_o <= x"05FD21D0";
      when 2225 => data_o <= x"7400004B";
      when 2226 => data_o <= x"052F400C";
      when 2227 => data_o <= x"D090DE20";
      when 2228 => data_o <= x"F4000200";
      when 2229 => data_o <= x"740000DA";
      when 2230 => data_o <= x"7400089A";
      when 2231 => data_o <= x"2BD0000A";
      when 2232 => data_o <= x"D090F6F6";
      when 2233 => data_o <= x"6E420000";
      when 2234 => data_o <= x"E95008DB";
      when 2235 => data_o <= x"7400065D";
      when 2236 => data_o <= x"E95008C4";
      when 2237 => data_o <= x"F3B74067";
      when 2238 => data_o <= x"444F4207";
      when 2239 => data_o <= x"203D2059";
      when 2240 => data_o <= x"39D0012C";
      when 2241 => data_o <= x"74000192";
      when 2242 => data_o <= x"74000148";
      when 2243 => data_o <= x"540008DB";
      when 2244 => data_o <= x"F1D00067";
      when 2245 => data_o <= x"20202015";
      when 2246 => data_o <= x"52432020";
      when 2247 => data_o <= x"45544145";
      when 2248 => data_o <= x"6C617620";
      when 2249 => data_o <= x"69206575";
      when 2250 => data_o <= x"FFFF2073";
      when 2251 => data_o <= x"39D0012C";
      when 2252 => data_o <= x"74000350";
      when 2253 => data_o <= x"B9D00192";
      when 2254 => data_o <= x"7400033E";
      when 2255 => data_o <= x"74000148";
      when 2256 => data_o <= x"74000067";
      when 2257 => data_o <= x"20202015";
      when 2258 => data_o <= x"4F442020";
      when 2259 => data_o <= x"203E5345";
      when 2260 => data_o <= x"69746361";
      when 2261 => data_o <= x"69206E6F";
      when 2262 => data_o <= x"FFFF3A73";
      when 2263 => data_o <= x"39D0012C";
      when 2264 => data_o <= x"74000148";
      when 2265 => data_o <= x"104F400A";
      when 2266 => data_o <= x"5400089A";
      when 2267 => data_o <= x"EC220000";
      when 2268 => data_o <= x"7400042C";
      when 2269 => data_o <= x"05FD09D0";
      when 2270 => data_o <= x"DBD00008";
      when 2271 => data_o <= x"7400009D";
      when 2272 => data_o <= x"4BD00005";
      when 2273 => data_o <= x"D090F60C";
      when 2274 => data_o <= x"74000067";
      when 2275 => data_o <= x"6E694C05";
      when 2276 => data_o <= x"FFFF2065";
      when 2277 => data_o <= x"39D0012C";
      when 2278 => data_o <= x"74000192";
      when 2279 => data_o <= x"2BD00009";
      when 2280 => data_o <= x"D090F620";
      when 2281 => data_o <= x"74000067";
      when 2282 => data_o <= x"6C694605";
      when 2283 => data_o <= x"FFFF2065";
      when 2284 => data_o <= x"39D0012C";
      when 2285 => data_o <= x"F4004000";
      when 2286 => data_o <= x"F3420000";
      when 2287 => data_o <= x"7EE28920";
      when 2288 => data_o <= x"C15008EF";
      when 2289 => data_o <= x"EE138800";
      when 2290 => data_o <= x"7400012C";
      when 2291 => data_o <= x"54000148";
      when 2292 => data_o <= x"F4000D9C";
      when 2293 => data_o <= x"D36F4000";
      when 2294 => data_o <= x"74000061";
      when 2295 => data_o <= x"540008FC";
      when 2296 => data_o <= x"F4009000";
      when 2297 => data_o <= x"74000594";
      when 2298 => data_o <= x"D090C800";
      when 2299 => data_o <= x"54000907";
      when 2300 => data_o <= x"F4000001";
      when 2301 => data_o <= x"74000061";
      when 2302 => data_o <= x"54000903";
      when 2303 => data_o <= x"F4004000";
      when 2304 => data_o <= x"74000594";
      when 2305 => data_o <= x"D090C800";
      when 2306 => data_o <= x"54000907";
      when 2307 => data_o <= x"F4000DE3";
      when 2308 => data_o <= x"D2EF8000";
      when 2309 => data_o <= x"D090FC20";
      when 2310 => data_o <= x"740004DE";
      when 2311 => data_o <= x"08800000";
      when 2312 => data_o <= x"04800000";
      when 2313 => data_o <= x"EBB08800";
      when 2314 => data_o <= x"F1FD09D0";
      when 2315 => data_o <= x"74000908";
      when 2316 => data_o <= x"2BC08800";
      when 2317 => data_o <= x"74000430";
      when 2318 => data_o <= x"5400030B";
      when 2319 => data_o <= x"04800000";
      when 2320 => data_o <= x"E9500914";
      when 2321 => data_o <= x"D09D39E7";
      when 2322 => data_o <= x"D9D00164";
      when 2323 => data_o <= x"5400090F";
      when 2324 => data_o <= x"EFB08800";
      when 2325 => data_o <= x"740003ED";
      when 2326 => data_o <= x"74000419";
      when 2327 => data_o <= x"EE408800";
      when 2328 => data_o <= x"74000915";
      when 2329 => data_o <= x"90220000";
      when 2330 => data_o <= x"7FC2BCF0";
      when 2331 => data_o <= x"E79740DD";
      when 2332 => data_o <= x"7F424328";
      when 2333 => data_o <= x"F1F7C800";
      when 2334 => data_o <= x"74000064";
      when 2335 => data_o <= x"54000928";
      when 2336 => data_o <= x"39FF0E7C";
      when 2337 => data_o <= x"F0A2B427";
      when 2338 => data_o <= x"04800000";
      when 2339 => data_o <= x"E9500927";
      when 2340 => data_o <= x"2BB2BB7C";
      when 2341 => data_o <= x"EFB2AC10";
      when 2342 => data_o <= x"24220000";
      when 2343 => data_o <= x"ED50091E";
      when 2344 => data_o <= x"EFB28120";
      when 2345 => data_o <= x"E950092B";
      when 2346 => data_o <= x"B0424220";
      when 2347 => data_o <= x"08800000";
      when 2348 => data_o <= x"F4000020";
      when 2349 => data_o <= x"5400008D";
      when 2350 => data_o <= x"E790F424";
      when 2351 => data_o <= x"D36F4020";
      when 2352 => data_o <= x"6E4E5320";
      when 2353 => data_o <= x"E9500934";
      when 2354 => data_o <= x"D09D0800";
      when 2355 => data_o <= x"5400092E";
      when 2356 => data_o <= x"08800000";
      when 2357 => data_o <= x"04800000";
      when 2358 => data_o <= x"EBB08800";
      when 2359 => data_o <= x"74000015";
      when 2360 => data_o <= x"E7920000";
      when 2361 => data_o <= x"04800000";
      when 2362 => data_o <= x"E9500949";
      when 2363 => data_o <= x"E7974019";
      when 2364 => data_o <= x"7FC2BCE4";
      when 2365 => data_o <= x"740000DA";
      when 2366 => data_o <= x"F1FF0A20";
      when 2367 => data_o <= x"7400091A";
      when 2368 => data_o <= x"90800000";
      when 2369 => data_o <= x"E9500946";
      when 2370 => data_o <= x"7400001D";
      when 2371 => data_o <= x"EFB74017";
      when 2372 => data_o <= x"EFBF4000";
      when 2373 => data_o <= x"D0220000";
      when 2374 => data_o <= x"F4000001";
      when 2375 => data_o <= x"740000E6";
      when 2376 => data_o <= x"54000939";
      when 2377 => data_o <= x"EFB74017";
      when 2378 => data_o <= x"EFBF4000";
      when 2379 => data_o <= x"08800000";
      when 2380 => data_o <= x"EC220000";
      when 2381 => data_o <= x"74000015";
      when 2382 => data_o <= x"7400001D";
      when 2383 => data_o <= x"74000017";
      when 2384 => data_o <= x"5400001D";
      when 2385 => data_o <= x"7400094D";
      when 2386 => data_o <= x"5400094D";
      when 2387 => data_o <= x"7400001D";
      when 2388 => data_o <= x"EFB08800";
      when 2389 => data_o <= x"7400001D";
      when 2390 => data_o <= x"5400001F";
      when 2391 => data_o <= x"74000035";
      when 2392 => data_o <= x"54000033";
      when 2393 => data_o <= x"74000957";
      when 2394 => data_o <= x"B0220000";
      when 2395 => data_o <= x"74000957";
      when 2396 => data_o <= x"90220000";
      when 2397 => data_o <= x"74000031";
      when 2398 => data_o <= x"90220000";
      when 2399 => data_o <= x"F3BB0220";
      when 2400 => data_o <= x"F04F0C08";
      when 2401 => data_o <= x"53C20000";
      when 2402 => data_o <= x"E1500964";
      when 2403 => data_o <= x"53C08800";
      when 2404 => data_o <= x"F4000080";
      when 2405 => data_o <= x"94000000";
      when 2406 => data_o <= x"74000031";
      when 2407 => data_o <= x"F0220000";
      when 2408 => data_o <= x"F1D005A8";
      when 2409 => data_o <= x"540005A8";
      when 2410 => data_o <= x"74000648";
      when 2411 => data_o <= x"F4000002";
      when 2412 => data_o <= x"10454598";
      when 2413 => data_o <= x"74000648";
      when 2414 => data_o <= x"74000270";
      when 2415 => data_o <= x"74000270";
      when 2416 => data_o <= x"74000668";
      when 2417 => data_o <= x"5400002D";
      when 2418 => data_o <= x"7FC2BCE4";
      when 2419 => data_o <= x"E5B90800";
      when 2420 => data_o <= x"E9500976";
      when 2421 => data_o <= x"EFB5406A";
      when 2422 => data_o <= x"74000953";
      when 2423 => data_o <= x"54000070";
      when 2424 => data_o <= x"7FC2BCE4";
      when 2425 => data_o <= x"E5B90800";
      when 2426 => data_o <= x"E950097C";
      when 2427 => data_o <= x"EFB5406A";
      when 2428 => data_o <= x"74000953";
      when 2429 => data_o <= x"F150006A";
      when 2430 => data_o <= x"7400001F";
      when 2431 => data_o <= x"7400001F";
      when 2432 => data_o <= x"74000972";
      when 2433 => data_o <= x"E9500983";
      when 2434 => data_o <= x"7400001D";
      when 2435 => data_o <= x"EFB08800";
      when 2436 => data_o <= x"7400001F";
      when 2437 => data_o <= x"7400001F";
      when 2438 => data_o <= x"74000972";
      when 2439 => data_o <= x"90800000";
      when 2440 => data_o <= x"E950098A";
      when 2441 => data_o <= x"7400001D";
      when 2442 => data_o <= x"EFB08800";
      when 2443 => data_o <= x"74000024";
      when 2444 => data_o <= x"54000033";
      when 2445 => data_o <= x"E796DF20";
      when 2446 => data_o <= x"7400002F";
      when 2447 => data_o <= x"F1D0002F";
      when 2448 => data_o <= x"740000A7";
      when 2449 => data_o <= x"2AC20000";
      when 2450 => data_o <= x"E9500994";
      when 2451 => data_o <= x"74000035";
      when 2452 => data_o <= x"08800000";
      when 2453 => data_o <= x"7F9E5D31";
      when 2454 => data_o <= x"04800000";
      when 2455 => data_o <= x"E950099A";
      when 2456 => data_o <= x"EDD00035";
      when 2457 => data_o <= x"F4000001";
      when 2458 => data_o <= x"283D0908";
      when 2459 => data_o <= x"E796DF7C";
      when 2460 => data_o <= x"74000038";
      when 2461 => data_o <= x"29D0002F";
      when 2462 => data_o <= x"74000015";
      when 2463 => data_o <= x"49D000A7";
      when 2464 => data_o <= x"F4000000";
      when 2465 => data_o <= x"74000017";
      when 2466 => data_o <= x"740000A7";
      when 2467 => data_o <= x"74000033";
      when 2468 => data_o <= x"2AC20000";
      when 2469 => data_o <= x"E95009A7";
      when 2470 => data_o <= x"74000995";
      when 2471 => data_o <= x"08800000";
      when 2472 => data_o <= x"E5F7C1B0";
      when 2473 => data_o <= x"E95009AB";
      when 2474 => data_o <= x"74000995";
      when 2475 => data_o <= x"49D000AC";
      when 2476 => data_o <= x"7FC2BC7C";
      when 2477 => data_o <= x"F0AF0A20";
      when 2478 => data_o <= x"740000AC";
      when 2479 => data_o <= x"F3BF0AB0";
      when 2480 => data_o <= x"E95009B2";
      when 2481 => data_o <= x"74000035";
      when 2482 => data_o <= x"08800000";
      when 2483 => data_o <= x"7DD0099B";
      when 2484 => data_o <= x"295009A8";
      when 2485 => data_o <= x"74000067";
      when 2486 => data_o <= x"79614D1A";
      when 2487 => data_o <= x"65687420";
      when 2488 => data_o <= x"726F4620";
      when 2489 => data_o <= x"62206874";
      when 2490 => data_o <= x"69772065";
      when 2491 => data_o <= x"79206874";
      when 2492 => data_o <= x"FF21756F";
      when 2493 => data_o <= x"39D0012C";
      when 2494 => data_o <= x"74000148";
      when 2495 => data_o <= x"5400072D";
      when 2496 => data_o <= x"07D00002";
      when 2497 => data_o <= x"74000070";
      when 2498 => data_o <= x"E95009C9";
      when 2499 => data_o <= x"07427420";
      when 2500 => data_o <= x"740009C0";
      when 2501 => data_o <= x"F3D00002";
      when 2502 => data_o <= x"D090C800";
      when 2503 => data_o <= x"740009C0";
      when 2504 => data_o <= x"0C220000";
      when 2505 => data_o <= x"EFD00001";
      when 2506 => data_o <= x"08800000";
      when 2507 => data_o <= x"F4000053";
      when 2508 => data_o <= x"94E2D623";
      when 2509 => data_o <= x"740000A7";
      when 2510 => data_o <= x"F3B08800";
      when 2511 => data_o <= x"74000116";
      when 2512 => data_o <= x"7FD0001E";
      when 2513 => data_o <= x"740009C0";
      when 2514 => data_o <= x"EDD00067";
      when 2515 => data_o <= x"20303313";
      when 2516 => data_o <= x"20626966";
      when 2517 => data_o <= x"63657865";
      when 2518 => data_o <= x"73657475";
      when 2519 => data_o <= x"206E6920";
      when 2520 => data_o <= x"39D0012C";
      when 2521 => data_o <= x"74000116";
      when 2522 => data_o <= x"2B424320";
      when 2523 => data_o <= x"740009CB";
      when 2524 => data_o <= x"F4000000";
      when 2525 => data_o <= x"74000161";
      when 2526 => data_o <= x"74000168";
      when 2527 => data_o <= x"F400002E";
      when 2528 => data_o <= x"74000164";
      when 2529 => data_o <= x"74000175";
      when 2530 => data_o <= x"7400017D";
      when 2531 => data_o <= x"7400012C";
      when 2532 => data_o <= x"74000067";
      when 2533 => data_o <= x"736D2006";
      when 2534 => data_o <= x"FF206365";
      when 2535 => data_o <= x"3950012C";
      when 2536 => data_o <= x"7FD00000";
      when 2537 => data_o <= x"F0800000";
      when 2538 => data_o <= x"10A31F80";
      when 2539 => data_o <= x"F0AF0220";
      when 2540 => data_o <= x"0416FC20";
      when 2541 => data_o <= x"120F0220";
      when 2542 => data_o <= x"00000003";
      when 2543 => data_o <= x"FFFFF204";
      when 2544 => data_o <= x"FFFFF200";
      when 2545 => data_o <= x"FFFFF1F0";
      when 2546 => data_o <= x"FFFFF100";
      when 2547 => data_o <= x"00000004";
      when 2548 => data_o <= x"FFFFF218";
      when 2549 => data_o <= x"0000000A";
      when 2550 => data_o <= x"000070B0";
      when 2551 => data_o <= x"000027DC";
      when 2552 => data_o <= x"FFFFF338";
      when 2553 => data_o <= x"00000006";
      when 2554 => data_o <= x"FFFFF22C";
      when 2555 => data_o <= x"FFFFF334";
      when 2556 => data_o <= x"000004F0";
      when 2557 => data_o <= x"00000001";
      when 2558 => data_o <= x"0000000C";
      when 2559 => data_o <= x"FFFFF26C";
      when 2560 => data_o <= x"0000000C";
      when 2561 => data_o <= x"00000001";
      when 2562 => data_o <= x"FFFFF248";
      when 2563 => data_o <= x"001A0001";
      when 2564 => data_o <= x"00000001";
      when 2565 => data_o <= x"FFFFF250";
      when 2566 => data_o <= x"140027A0";
      when 2567 => data_o <= x"00000003";
      when 2568 => data_o <= x"FFFFF25C";
      when 2569 => data_o <= x"000055E8";
      when 2570 => data_o <= x"00140003";
      when 2571 => data_o <= x"FFFFF334";
      when 2572 => data_o <= x"00000001";
      when 2573 => data_o <= x"FFFFF334";
      when 2574 => data_o <= x"00007090";
      when 2575 => data_o <= x"00000000";
      when 2576 => data_o <= x"FFFFF338";
      when 2577 => data_o <= x"F4000DFF";
      when 2578 => data_o <= x"D01D0920";
      when 2579 => data_o <= x"74000093";
      when 2580 => data_o <= x"F40027B8";
      when 2581 => data_o <= x"9B9E4910";
      when 2582 => data_o <= x"103F1FF0";
      when 2583 => data_o <= x"28120000";
      when 2584 => data_o <= x"E9500A1B";
      when 2585 => data_o <= x"7E629D71";
      when 2586 => data_o <= x"54000A15";
      when 2587 => data_o <= x"2BD00D97";
      when 2588 => data_o <= x"D27EC800";
      when 2589 => data_o <= x"F4000DFF";
      when 2590 => data_o <= x"D3FF4EFF";
      when 2591 => data_o <= x"D37F4E13";
      when 2592 => data_o <= x"D2FF4D97";
      when 2593 => data_o <= x"D2E7C800";
      when 2594 => data_o <= x"F4010000";
      when 2595 => data_o <= x"F4000DDF";
      when 2596 => data_o <= x"D27EC800";
      when 2597 => data_o <= x"F4018000";
      when 2598 => data_o <= x"F4000DE3";
      when 2599 => data_o <= x"D27EC220";
      when 2600 => data_o <= x"74000A11";
      when 2601 => data_o <= x"740009B5";
      when 2602 => data_o <= x"540000F6";
      when 2603 => data_o <= x"74000A11";
      when 2604 => data_o <= x"740009B5";
      when 2605 => data_o <= x"540000F6";
      when 2606 => data_o <= x"FFFFFFFF";
      when 2607 => data_o <= x"FFFFFFFF";
      when 2608 => data_o <= x"FFFFFFFF";
      when 2609 => data_o <= x"FFFFFFFF";
      when 2610 => data_o <= x"FFFFFFFF";
      when 2611 => data_o <= x"FFFFFFFF";
      when 2612 => data_o <= x"FFFFFFFF";
      when 2613 => data_o <= x"FFFFFFFF";
      when 2614 => data_o <= x"FFFFFFFF";
      when 2615 => data_o <= x"FFFFFFFF";
      when 2616 => data_o <= x"FFFFFFFF";
      when 2617 => data_o <= x"FFFFFFFF";
      when 2618 => data_o <= x"FFFFFFFF";
      when 2619 => data_o <= x"FFFFFFFF";
      when 2620 => data_o <= x"FFFFFFFF";
      when 2621 => data_o <= x"FFFFFFFF";
      when 2622 => data_o <= x"FFFFFFFF";
      when 2623 => data_o <= x"FFFFFFFF";
      when 2624 => data_o <= x"FFFFFFFF";
      when 2625 => data_o <= x"FFFFFFFF";
      when 2626 => data_o <= x"FFFFFFFF";
      when 2627 => data_o <= x"FFFFFFFF";
      when 2628 => data_o <= x"FFFFFFFF";
      when 2629 => data_o <= x"FFFFFFFF";
      when 2630 => data_o <= x"FFFFFFFF";
      when 2631 => data_o <= x"FFFFFFFF";
      when 2632 => data_o <= x"FFFFFFFF";
      when 2633 => data_o <= x"FFFFFFFF";
      when 2634 => data_o <= x"FFFFFFFF";
      when 2635 => data_o <= x"FFFFFFFF";
      when 2636 => data_o <= x"FFFFFFFF";
      when 2637 => data_o <= x"FFFFFFFF";
      when 2638 => data_o <= x"FFFFFFFF";
      when 2639 => data_o <= x"FFFFFFFF";
      when 2640 => data_o <= x"FFFFFFFF";
      when 2641 => data_o <= x"FFFFFFFF";
      when 2642 => data_o <= x"FFFFFFFF";
      when 2643 => data_o <= x"FFFFFFFF";
      when 2644 => data_o <= x"FFFFFFFF";
      when 2645 => data_o <= x"FFFFFFFF";
      when 2646 => data_o <= x"FFFFFFFF";
      when 2647 => data_o <= x"FFFFFFFF";
      when 2648 => data_o <= x"FFFFFFFF";
      when 2649 => data_o <= x"FFFFFFFF";
      when 2650 => data_o <= x"FFFFFFFF";
      when 2651 => data_o <= x"FFFFFFFF";
      when 2652 => data_o <= x"FFFFFFFF";
      when 2653 => data_o <= x"FFFFFFFF";
      when 2654 => data_o <= x"FFFFFFFF";
      when 2655 => data_o <= x"FFFFFFFF";
      when 2656 => data_o <= x"FFFFFFFF";
      when 2657 => data_o <= x"FFFFFFFF";
      when 2658 => data_o <= x"FFFFFFFF";
      when 2659 => data_o <= x"FFFFFFFF";
      when 2660 => data_o <= x"FFFFFFFF";
      when 2661 => data_o <= x"FFFFFFFF";
      when 2662 => data_o <= x"FFFFFFFF";
      when 2663 => data_o <= x"FFFFFFFF";
      when 2664 => data_o <= x"FFFFFFFF";
      when 2665 => data_o <= x"FFFFFFFF";
      when 2666 => data_o <= x"FFFFFFFF";
      when 2667 => data_o <= x"FFFFFFFF";
      when 2668 => data_o <= x"FFFFFFFF";
      when 2669 => data_o <= x"FFFFFFFF";
      when 2670 => data_o <= x"FFFFFFFF";
      when 2671 => data_o <= x"FFFFFFFF";
      when 2672 => data_o <= x"FFFFFFFF";
      when 2673 => data_o <= x"FFFFFFFF";
      when 2674 => data_o <= x"FFFFFFFF";
      when 2675 => data_o <= x"FFFFFFFF";
      when 2676 => data_o <= x"FFFFFFFF";
      when 2677 => data_o <= x"FFFFFFFF";
      when 2678 => data_o <= x"FFFFFFFF";
      when 2679 => data_o <= x"FFFFFFFF";
      when 2680 => data_o <= x"FFFFFFFF";
      when 2681 => data_o <= x"FFFFFFFF";
      when 2682 => data_o <= x"FFFFFFFF";
      when 2683 => data_o <= x"FFFFFFFF";
      when 2684 => data_o <= x"FFFFFFFF";
      when 2685 => data_o <= x"FFFFFFFF";
      when 2686 => data_o <= x"FFFFFFFF";
      when 2687 => data_o <= x"FFFFFFFF";
      when 2688 => data_o <= x"FFFFFFFF";
      when 2689 => data_o <= x"FFFFFFFF";
      when 2690 => data_o <= x"FFFFFFFF";
      when 2691 => data_o <= x"FFFFFFFF";
      when 2692 => data_o <= x"FFFFFFFF";
      when 2693 => data_o <= x"FFFFFFFF";
      when 2694 => data_o <= x"FFFFFFFF";
      when 2695 => data_o <= x"FFFFFFFF";
      when 2696 => data_o <= x"FFFFFFFF";
      when 2697 => data_o <= x"FFFFFFFF";
      when 2698 => data_o <= x"FFFFFFFF";
      when 2699 => data_o <= x"FFFFFFFF";
      when 2700 => data_o <= x"FFFFFFFF";
      when 2701 => data_o <= x"FFFFFFFF";
      when 2702 => data_o <= x"FFFFFFFF";
      when 2703 => data_o <= x"FFFFFFFF";
      when 2704 => data_o <= x"FFFFFFFF";
      when 2705 => data_o <= x"FFFFFFFF";
      when 2706 => data_o <= x"FFFFFFFF";
      when 2707 => data_o <= x"FFFFFFFF";
      when 2708 => data_o <= x"FFFFFFFF";
      when 2709 => data_o <= x"FFFFFFFF";
      when 2710 => data_o <= x"FFFFFFFF";
      when 2711 => data_o <= x"FFFFFFFF";
      when 2712 => data_o <= x"FFFFFFFF";
      when 2713 => data_o <= x"FFFFFFFF";
      when 2714 => data_o <= x"FFFFFFFF";
      when 2715 => data_o <= x"FFFFFFFF";
      when 2716 => data_o <= x"FFFFFFFF";
      when 2717 => data_o <= x"FFFFFFFF";
      when 2718 => data_o <= x"FFFFFFFF";
      when 2719 => data_o <= x"FFFFFFFF";
      when 2720 => data_o <= x"FFFFFFFF";
      when 2721 => data_o <= x"FFFFFFFF";
      when 2722 => data_o <= x"FFFFFFFF";
      when 2723 => data_o <= x"FFFFFFFF";
      when 2724 => data_o <= x"FFFFFFFF";
      when 2725 => data_o <= x"FFFFFFFF";
      when 2726 => data_o <= x"FFFFFFFF";
      when 2727 => data_o <= x"FFFFFFFF";
      when 2728 => data_o <= x"FFFFFFFF";
      when 2729 => data_o <= x"FFFFFFFF";
      when 2730 => data_o <= x"FFFFFFFF";
      when 2731 => data_o <= x"FFFFFFFF";
      when 2732 => data_o <= x"FFFFFFFF";
      when 2733 => data_o <= x"FFFFFFFF";
      when 2734 => data_o <= x"FFFFFFFF";
      when 2735 => data_o <= x"FFFFFFFF";
      when 2736 => data_o <= x"FFFFFFFF";
      when 2737 => data_o <= x"FFFFFFFF";
      when 2738 => data_o <= x"FFFFFFFF";
      when 2739 => data_o <= x"FFFFFFFF";
      when 2740 => data_o <= x"FFFFFFFF";
      when 2741 => data_o <= x"FFFFFFFF";
      when 2742 => data_o <= x"FFFFFFFF";
      when 2743 => data_o <= x"FFFFFFFF";
      when 2744 => data_o <= x"FFFFFFFF";
      when 2745 => data_o <= x"FFFFFFFF";
      when 2746 => data_o <= x"FFFFFFFF";
      when 2747 => data_o <= x"FFFFFFFF";
      when 2748 => data_o <= x"FFFFFFFF";
      when 2749 => data_o <= x"FFFFFFFF";
      when 2750 => data_o <= x"FFFFFFFF";
      when 2751 => data_o <= x"FFFFFFFF";
      when 2752 => data_o <= x"FFFFFFFF";
      when 2753 => data_o <= x"FFFFFFFF";
      when 2754 => data_o <= x"FFFFFFFF";
      when 2755 => data_o <= x"FFFFFFFF";
      when 2756 => data_o <= x"FFFFFFFF";
      when 2757 => data_o <= x"FFFFFFFF";
      when 2758 => data_o <= x"FFFFFFFF";
      when 2759 => data_o <= x"FFFFFFFF";
      when 2760 => data_o <= x"FFFFFFFF";
      when 2761 => data_o <= x"FFFFFFFF";
      when 2762 => data_o <= x"FFFFFFFF";
      when 2763 => data_o <= x"FFFFFFFF";
      when 2764 => data_o <= x"FFFFFFFF";
      when 2765 => data_o <= x"FFFFFFFF";
      when 2766 => data_o <= x"FFFFFFFF";
      when 2767 => data_o <= x"FFFFFFFF";
      when 2768 => data_o <= x"FFFFFFFF";
      when 2769 => data_o <= x"FFFFFFFF";
      when 2770 => data_o <= x"FFFFFFFF";
      when 2771 => data_o <= x"FFFFFFFF";
      when 2772 => data_o <= x"FFFFFFFF";
      when 2773 => data_o <= x"FFFFFFFF";
      when 2774 => data_o <= x"FFFFFFFF";
      when 2775 => data_o <= x"FFFFFFFF";
      when 2776 => data_o <= x"FFFFFFFF";
      when 2777 => data_o <= x"FFFFFFFF";
      when 2778 => data_o <= x"FFFFFFFF";
      when 2779 => data_o <= x"FFFFFFFF";
      when 2780 => data_o <= x"FFFFFFFF";
      when 2781 => data_o <= x"FFFFFFFF";
      when 2782 => data_o <= x"FFFFFFFF";
      when 2783 => data_o <= x"FFFFFFFF";
      when 2784 => data_o <= x"FFFFFFFF";
      when 2785 => data_o <= x"FFFFFFFF";
      when 2786 => data_o <= x"FFFFFFFF";
      when 2787 => data_o <= x"FFFFFFFF";
      when 2788 => data_o <= x"FFFFFFFF";
      when 2789 => data_o <= x"FFFFFFFF";
      when 2790 => data_o <= x"FFFFFFFF";
      when 2791 => data_o <= x"FFFFFFFF";
      when 2792 => data_o <= x"FFFFFFFF";
      when 2793 => data_o <= x"FFFFFFFF";
      when 2794 => data_o <= x"FFFFFFFF";
      when 2795 => data_o <= x"FFFFFFFF";
      when 2796 => data_o <= x"FFFFFFFF";
      when 2797 => data_o <= x"FFFFFFFF";
      when 2798 => data_o <= x"FFFFFFFF";
      when 2799 => data_o <= x"FFFFFFFF";
      when 2800 => data_o <= x"FFFFFFFF";
      when 2801 => data_o <= x"FFFFFFFF";
      when 2802 => data_o <= x"FFFFFFFF";
      when 2803 => data_o <= x"FFFFFFFF";
      when 2804 => data_o <= x"FFFFFFFF";
      when 2805 => data_o <= x"FFFFFFFF";
      when 2806 => data_o <= x"FFFFFFFF";
      when 2807 => data_o <= x"FFFFFFFF";
      when 2808 => data_o <= x"FFFFFFFF";
      when 2809 => data_o <= x"FFFFFFFF";
      when 2810 => data_o <= x"FFFFFFFF";
      when 2811 => data_o <= x"FFFFFFFF";
      when 2812 => data_o <= x"FFFFFFFF";
      when 2813 => data_o <= x"FFFFFFFF";
      when 2814 => data_o <= x"FFFFFFFF";
      when 2815 => data_o <= x"FFFFFFFF";
      when 2816 => data_o <= x"FFFFFFFF";
      when 2817 => data_o <= x"FFFFFFFF";
      when 2818 => data_o <= x"FFFFFFFF";
      when 2819 => data_o <= x"FFFFFFFF";
      when 2820 => data_o <= x"FFFFFFFF";
      when 2821 => data_o <= x"FFFFFFFF";
      when 2822 => data_o <= x"FFFFFFFF";
      when 2823 => data_o <= x"FFFFFFFF";
      when 2824 => data_o <= x"FFFFFFFF";
      when 2825 => data_o <= x"FFFFFFFF";
      when 2826 => data_o <= x"FFFFFFFF";
      when 2827 => data_o <= x"FFFFFFFF";
      when 2828 => data_o <= x"FFFFFFFF";
      when 2829 => data_o <= x"FFFFFFFF";
      when 2830 => data_o <= x"FFFFFFFF";
      when 2831 => data_o <= x"FFFFFFFF";
      when 2832 => data_o <= x"FFFFFFFF";
      when 2833 => data_o <= x"FFFFFFFF";
      when 2834 => data_o <= x"FFFFFFFF";
      when 2835 => data_o <= x"FFFFFFFF";
      when 2836 => data_o <= x"FFFFFFFF";
      when 2837 => data_o <= x"FFFFFFFF";
      when 2838 => data_o <= x"FFFFFFFF";
      when 2839 => data_o <= x"FFFFFFFF";
      when 2840 => data_o <= x"FFFFFFFF";
      when 2841 => data_o <= x"FFFFFFFF";
      when 2842 => data_o <= x"FFFFFFFF";
      when 2843 => data_o <= x"FFFFFFFF";
      when 2844 => data_o <= x"FFFFFFFF";
      when 2845 => data_o <= x"FFFFFFFF";
      when 2846 => data_o <= x"FFFFFFFF";
      when 2847 => data_o <= x"FFFFFFFF";
      when 2848 => data_o <= x"FFFFFFFF";
      when 2849 => data_o <= x"FFFFFFFF";
      when 2850 => data_o <= x"FFFFFFFF";
      when 2851 => data_o <= x"FFFFFFFF";
      when 2852 => data_o <= x"FFFFFFFF";
      when 2853 => data_o <= x"FFFFFFFF";
      when 2854 => data_o <= x"FFFFFFFF";
      when 2855 => data_o <= x"FFFFFFFF";
      when 2856 => data_o <= x"FFFFFFFF";
      when 2857 => data_o <= x"FFFFFFFF";
      when 2858 => data_o <= x"FFFFFFFF";
      when 2859 => data_o <= x"FFFFFFFF";
      when 2860 => data_o <= x"FFFFFFFF";
      when 2861 => data_o <= x"FFFFFFFF";
      when 2862 => data_o <= x"FFFFFFFF";
      when 2863 => data_o <= x"FFFFFFFF";
      when 2864 => data_o <= x"FFFFFFFF";
      when 2865 => data_o <= x"FFFFFFFF";
      when 2866 => data_o <= x"FFFFFFFF";
      when 2867 => data_o <= x"FFFFFFFF";
      when 2868 => data_o <= x"FFFFFFFF";
      when 2869 => data_o <= x"FFFFFFFF";
      when 2870 => data_o <= x"FFFFFFFF";
      when 2871 => data_o <= x"FFFFFFFF";
      when 2872 => data_o <= x"FFFFFFFF";
      when 2873 => data_o <= x"FFFFFFFF";
      when 2874 => data_o <= x"FFFFFFFF";
      when 2875 => data_o <= x"FFFFFFFF";
      when 2876 => data_o <= x"FFFFFFFF";
      when 2877 => data_o <= x"FFFFFFFF";
      when 2878 => data_o <= x"FFFFFFFF";
      when 2879 => data_o <= x"FFFFFFFF";
      when 2880 => data_o <= x"FFFFFFFF";
      when 2881 => data_o <= x"FFFFFFFF";
      when 2882 => data_o <= x"FFFFFFFF";
      when 2883 => data_o <= x"FFFFFFFF";
      when 2884 => data_o <= x"FFFFFFFF";
      when 2885 => data_o <= x"FFFFFFFF";
      when 2886 => data_o <= x"FFFFFFFF";
      when 2887 => data_o <= x"FFFFFFFF";
      when 2888 => data_o <= x"FFFFFFFF";
      when 2889 => data_o <= x"FFFFFFFF";
      when 2890 => data_o <= x"FFFFFFFF";
      when 2891 => data_o <= x"FFFFFFFF";
      when 2892 => data_o <= x"FFFFFFFF";
      when 2893 => data_o <= x"FFFFFFFF";
      when 2894 => data_o <= x"FFFFFFFF";
      when 2895 => data_o <= x"FFFFFFFF";
      when 2896 => data_o <= x"FFFFFFFF";
      when 2897 => data_o <= x"FFFFFFFF";
      when 2898 => data_o <= x"FFFFFFFF";
      when 2899 => data_o <= x"FFFFFFFF";
      when 2900 => data_o <= x"FFFFFFFF";
      when 2901 => data_o <= x"FFFFFFFF";
      when 2902 => data_o <= x"FFFFFFFF";
      when 2903 => data_o <= x"FFFFFFFF";
      when 2904 => data_o <= x"FFFFFFFF";
      when 2905 => data_o <= x"FFFFFFFF";
      when 2906 => data_o <= x"FFFFFFFF";
      when 2907 => data_o <= x"FFFFFFFF";
      when 2908 => data_o <= x"FFFFFFFF";
      when 2909 => data_o <= x"FFFFFFFF";
      when 2910 => data_o <= x"FFFFFFFF";
      when 2911 => data_o <= x"FFFFFFFF";
      when 2912 => data_o <= x"FFFFFFFF";
      when 2913 => data_o <= x"FFFFFFFF";
      when 2914 => data_o <= x"FFFFFFFF";
      when 2915 => data_o <= x"FFFFFFFF";
      when 2916 => data_o <= x"FFFFFFFF";
      when 2917 => data_o <= x"FFFFFFFF";
      when 2918 => data_o <= x"FFFFFFFF";
      when 2919 => data_o <= x"FFFFFFFF";
      when 2920 => data_o <= x"FFFFFFFF";
      when 2921 => data_o <= x"FFFFFFFF";
      when 2922 => data_o <= x"FFFFFFFF";
      when 2923 => data_o <= x"FFFFFFFF";
      when 2924 => data_o <= x"FFFFFFFF";
      when 2925 => data_o <= x"FFFFFFFF";
      when 2926 => data_o <= x"FFFFFFFF";
      when 2927 => data_o <= x"FFFFFFFF";
      when 2928 => data_o <= x"FFFFFFFF";
      when 2929 => data_o <= x"FFFFFFFF";
      when 2930 => data_o <= x"FFFFFFFF";
      when 2931 => data_o <= x"FFFFFFFF";
      when 2932 => data_o <= x"FFFFFFFF";
      when 2933 => data_o <= x"FFFFFFFF";
      when 2934 => data_o <= x"FFFFFFFF";
      when 2935 => data_o <= x"FFFFFFFF";
      when 2936 => data_o <= x"FFFFFFFF";
      when 2937 => data_o <= x"FFFFFFFF";
      when 2938 => data_o <= x"FFFFFFFF";
      when 2939 => data_o <= x"FFFFFFFF";
      when 2940 => data_o <= x"FFFFFFFF";
      when 2941 => data_o <= x"FFFFFFFF";
      when 2942 => data_o <= x"FFFFFFFF";
      when 2943 => data_o <= x"FFFFFFFF";
      when 2944 => data_o <= x"FFFFFFFF";
      when 2945 => data_o <= x"FFFFFFFF";
      when 2946 => data_o <= x"FFFFFFFF";
      when 2947 => data_o <= x"FFFFFFFF";
      when 2948 => data_o <= x"FFFFFFFF";
      when 2949 => data_o <= x"FFFFFFFF";
      when 2950 => data_o <= x"FFFFFFFF";
      when 2951 => data_o <= x"FFFFFFFF";
      when 2952 => data_o <= x"FFFFFFFF";
      when 2953 => data_o <= x"FFFFFFFF";
      when 2954 => data_o <= x"FFFFFFFF";
      when 2955 => data_o <= x"FFFFFFFF";
      when 2956 => data_o <= x"FFFFFFFF";
      when 2957 => data_o <= x"FFFFFFFF";
      when 2958 => data_o <= x"FFFFFFFF";
      when 2959 => data_o <= x"FFFFFFFF";
      when 2960 => data_o <= x"FFFFFFFF";
      when 2961 => data_o <= x"FFFFFFFF";
      when 2962 => data_o <= x"FFFFFFFF";
      when 2963 => data_o <= x"FFFFFFFF";
      when 2964 => data_o <= x"FFFFFFFF";
      when 2965 => data_o <= x"FFFFFFFF";
      when 2966 => data_o <= x"FFFFFFFF";
      when 2967 => data_o <= x"FFFFFFFF";
      when 2968 => data_o <= x"FFFFFFFF";
      when 2969 => data_o <= x"FFFFFFFF";
      when 2970 => data_o <= x"FFFFFFFF";
      when 2971 => data_o <= x"FFFFFFFF";
      when 2972 => data_o <= x"FFFFFFFF";
      when 2973 => data_o <= x"FFFFFFFF";
      when 2974 => data_o <= x"FFFFFFFF";
      when 2975 => data_o <= x"FFFFFFFF";
      when 2976 => data_o <= x"FFFFFFFF";
      when 2977 => data_o <= x"FFFFFFFF";
      when 2978 => data_o <= x"FFFFFFFF";
      when 2979 => data_o <= x"FFFFFFFF";
      when 2980 => data_o <= x"FFFFFFFF";
      when 2981 => data_o <= x"FFFFFFFF";
      when 2982 => data_o <= x"FFFFFFFF";
      when 2983 => data_o <= x"FFFFFFFF";
      when 2984 => data_o <= x"FFFFFFFF";
      when 2985 => data_o <= x"FFFFFFFF";
      when 2986 => data_o <= x"FFFFFFFF";
      when 2987 => data_o <= x"FFFFFFFF";
      when 2988 => data_o <= x"FFFFFFFF";
      when 2989 => data_o <= x"FFFFFFFF";
      when 2990 => data_o <= x"FFFFFFFF";
      when 2991 => data_o <= x"FFFFFFFF";
      when 2992 => data_o <= x"FFFFFFFF";
      when 2993 => data_o <= x"FFFFFFFF";
      when 2994 => data_o <= x"FFFFFFFF";
      when 2995 => data_o <= x"FFFFFFFF";
      when 2996 => data_o <= x"FFFFFFFF";
      when 2997 => data_o <= x"FFFFFFFF";
      when 2998 => data_o <= x"FFFFFFFF";
      when 2999 => data_o <= x"FFFFFFFF";
      when 3000 => data_o <= x"FFFFFFFF";
      when 3001 => data_o <= x"FFFFFFFF";
      when 3002 => data_o <= x"FFFFFFFF";
      when 3003 => data_o <= x"FFFFFFFF";
      when 3004 => data_o <= x"FFFFFFFF";
      when 3005 => data_o <= x"FFFFFFFF";
      when 3006 => data_o <= x"FFFFFFFF";
      when 3007 => data_o <= x"FFFFFFFF";
      when 3008 => data_o <= x"FFFFFFFF";
      when 3009 => data_o <= x"FFFFFFFF";
      when 3010 => data_o <= x"FFFFFFFF";
      when 3011 => data_o <= x"FFFFFFFF";
      when 3012 => data_o <= x"FFFFFFFF";
      when 3013 => data_o <= x"FFFFFFFF";
      when 3014 => data_o <= x"FFFFFFFF";
      when 3015 => data_o <= x"FFFFFFFF";
      when 3016 => data_o <= x"FFFFFFFF";
      when 3017 => data_o <= x"FFFFFFFF";
      when 3018 => data_o <= x"FFFFFFFF";
      when 3019 => data_o <= x"FFFFFFFF";
      when 3020 => data_o <= x"FFFFFFFF";
      when 3021 => data_o <= x"FFFFFFFF";
      when 3022 => data_o <= x"FFFFFFFF";
      when 3023 => data_o <= x"FFFFFFFF";
      when 3024 => data_o <= x"FFFFFFFF";
      when 3025 => data_o <= x"FFFFFFFF";
      when 3026 => data_o <= x"FFFFFFFF";
      when 3027 => data_o <= x"FFFFFFFF";
      when 3028 => data_o <= x"FFFFFFFF";
      when 3029 => data_o <= x"FFFFFFFF";
      when 3030 => data_o <= x"FFFFFFFF";
      when 3031 => data_o <= x"FFFFFFFF";
      when 3032 => data_o <= x"FFFFFFFF";
      when 3033 => data_o <= x"FFFFFFFF";
      when 3034 => data_o <= x"FFFFFFFF";
      when 3035 => data_o <= x"FFFFFFFF";
      when 3036 => data_o <= x"FFFFFFFF";
      when 3037 => data_o <= x"FFFFFFFF";
      when 3038 => data_o <= x"FFFFFFFF";
      when 3039 => data_o <= x"FFFFFFFF";
      when 3040 => data_o <= x"FFFFFFFF";
      when 3041 => data_o <= x"FFFFFFFF";
      when 3042 => data_o <= x"FFFFFFFF";
      when 3043 => data_o <= x"FFFFFFFF";
      when 3044 => data_o <= x"FFFFFFFF";
      when 3045 => data_o <= x"FFFFFFFF";
      when 3046 => data_o <= x"FFFFFFFF";
      when 3047 => data_o <= x"FFFFFFFF";
      when 3048 => data_o <= x"FFFFFFFF";
      when 3049 => data_o <= x"FFFFFFFF";
      when 3050 => data_o <= x"FFFFFFFF";
      when 3051 => data_o <= x"FFFFFFFF";
      when 3052 => data_o <= x"FFFFFFFF";
      when 3053 => data_o <= x"FFFFFFFF";
      when 3054 => data_o <= x"FFFFFFFF";
      when 3055 => data_o <= x"FFFFFFFF";
      when 3056 => data_o <= x"FFFFFFFF";
      when 3057 => data_o <= x"FFFFFFFF";
      when 3058 => data_o <= x"FFFFFFFF";
      when 3059 => data_o <= x"FFFFFFFF";
      when 3060 => data_o <= x"FFFFFFFF";
      when 3061 => data_o <= x"FFFFFFFF";
      when 3062 => data_o <= x"FFFFFFFF";
      when 3063 => data_o <= x"FFFFFFFF";
      when 3064 => data_o <= x"FFFFFFFF";
      when 3065 => data_o <= x"FFFFFFFF";
      when 3066 => data_o <= x"FFFFFFFF";
      when 3067 => data_o <= x"FFFFFFFF";
      when 3068 => data_o <= x"FFFFFFFF";
      when 3069 => data_o <= x"FFFFFFFF";
      when 3070 => data_o <= x"FFFFFFFF";
      when 3071 => data_o <= x"FFFFFFFF";
      when 3072 => data_o <= x"FFFFFFFF";
      when 3073 => data_o <= x"FFFFFFFF";
      when 3074 => data_o <= x"FFFFFFFF";
      when 3075 => data_o <= x"FFFFFFFF";
      when 3076 => data_o <= x"FFFFFFFF";
      when 3077 => data_o <= x"FFFFFFFF";
      when 3078 => data_o <= x"FFFFFFFF";
      when 3079 => data_o <= x"FFFFFFFF";
      when 3080 => data_o <= x"FFFFFFFF";
      when 3081 => data_o <= x"FFFFFFFF";
      when 3082 => data_o <= x"FFFFFFFF";
      when 3083 => data_o <= x"FFFFFFFF";
      when 3084 => data_o <= x"FFFFFFFF";
      when 3085 => data_o <= x"FFFFFFFF";
      when 3086 => data_o <= x"FFFFFFFF";
      when 3087 => data_o <= x"FFFFFFFF";
      when 3088 => data_o <= x"FFFFFFFF";
      when 3089 => data_o <= x"FFFFFFFF";
      when 3090 => data_o <= x"FFFFFFFF";
      when 3091 => data_o <= x"FFFFFFFF";
      when 3092 => data_o <= x"FFFFFFFF";
      when 3093 => data_o <= x"FFFFFFFF";
      when 3094 => data_o <= x"FFFFFFFF";
      when 3095 => data_o <= x"FFFFFFFF";
      when 3096 => data_o <= x"FFFFFFFF";
      when 3097 => data_o <= x"FFFFFFFF";
      when 3098 => data_o <= x"FFFFFFFF";
      when 3099 => data_o <= x"FFFFFFFF";
      when 3100 => data_o <= x"FFFFFFFF";
      when 3101 => data_o <= x"FFFFFFFF";
      when 3102 => data_o <= x"FFFFFFFF";
      when 3103 => data_o <= x"FFFFFFFF";
      when 3104 => data_o <= x"FFFFFFFF";
      when 3105 => data_o <= x"FFFFFFFF";
      when 3106 => data_o <= x"FFFFFFFF";
      when 3107 => data_o <= x"FFFFFFFF";
      when 3108 => data_o <= x"FFFFFFFF";
      when 3109 => data_o <= x"FFFFFFFF";
      when 3110 => data_o <= x"FFFFFFFF";
      when 3111 => data_o <= x"FFFFFFFF";
      when 3112 => data_o <= x"FFFFFFFF";
      when 3113 => data_o <= x"FFFFFFFF";
      when 3114 => data_o <= x"FFFFFFFF";
      when 3115 => data_o <= x"FFFFFFFF";
      when 3116 => data_o <= x"FFFFFFFF";
      when 3117 => data_o <= x"FFFFFFFF";
      when 3118 => data_o <= x"FFFFFFFF";
      when 3119 => data_o <= x"FFFFFFFF";
      when 3120 => data_o <= x"FFFFFFFF";
      when 3121 => data_o <= x"FFFFFFFF";
      when 3122 => data_o <= x"FFFFFFFF";
      when 3123 => data_o <= x"FFFFFFFF";
      when 3124 => data_o <= x"FFFFFFFF";
      when 3125 => data_o <= x"FFFFFFFF";
      when 3126 => data_o <= x"FFFFFFFF";
      when 3127 => data_o <= x"FFFFFFFF";
      when 3128 => data_o <= x"FFFFFFFF";
      when 3129 => data_o <= x"FFFFFFFF";
      when 3130 => data_o <= x"FFFFFFFF";
      when 3131 => data_o <= x"FFFFFFFF";
      when 3132 => data_o <= x"FFFFFFFF";
      when 3133 => data_o <= x"FFFFFFFF";
      when 3134 => data_o <= x"FFFFFFFF";
      when 3135 => data_o <= x"FFFFFFFF";
      when 3136 => data_o <= x"FFFFFFFF";
      when 3137 => data_o <= x"FFFFFFFF";
      when 3138 => data_o <= x"FFFFFFFF";
      when 3139 => data_o <= x"FFFFFFFF";
      when 3140 => data_o <= x"FFFFFFFF";
      when 3141 => data_o <= x"FFFFFFFF";
      when 3142 => data_o <= x"FFFFFFFF";
      when 3143 => data_o <= x"FFFFFFFF";
      when 3144 => data_o <= x"FFFFFFFF";
      when 3145 => data_o <= x"FFFFFFFF";
      when 3146 => data_o <= x"FFFFFFFF";
      when 3147 => data_o <= x"FFFFFFFF";
      when 3148 => data_o <= x"FFFFFFFF";
      when 3149 => data_o <= x"FFFFFFFF";
      when 3150 => data_o <= x"FFFFFFFF";
      when 3151 => data_o <= x"FFFFFFFF";
      when 3152 => data_o <= x"FFFFFFFF";
      when 3153 => data_o <= x"FFFFFFFF";
      when 3154 => data_o <= x"FFFFFFFF";
      when 3155 => data_o <= x"FFFFFFFF";
      when 3156 => data_o <= x"FFFFFFFF";
      when 3157 => data_o <= x"FFFFFFFF";
      when 3158 => data_o <= x"FFFFFFFF";
      when 3159 => data_o <= x"FFFFFFFF";
      when 3160 => data_o <= x"FFFFFFFF";
      when 3161 => data_o <= x"FFFFFFFF";
      when 3162 => data_o <= x"FFFFFFFF";
      when 3163 => data_o <= x"FFFFFFFF";
      when 3164 => data_o <= x"FFFFFFFF";
      when 3165 => data_o <= x"FFFFFFFF";
      when 3166 => data_o <= x"FFFFFFFF";
      when 3167 => data_o <= x"FFFFFFFF";
      when 3168 => data_o <= x"FFFFFFFF";
      when 3169 => data_o <= x"FFFFFFFF";
      when 3170 => data_o <= x"FFFFFFFF";
      when 3171 => data_o <= x"FFFFFFFF";
      when 3172 => data_o <= x"FFFFFFFF";
      when 3173 => data_o <= x"FFFFFFFF";
      when 3174 => data_o <= x"FFFFFFFF";
      when 3175 => data_o <= x"FFFFFFFF";
      when 3176 => data_o <= x"FFFFFFFF";
      when 3177 => data_o <= x"FFFFFFFF";
      when 3178 => data_o <= x"FFFFFFFF";
      when 3179 => data_o <= x"FFFFFFFF";
      when 3180 => data_o <= x"FFFFFFFF";
      when 3181 => data_o <= x"FFFFFFFF";
      when 3182 => data_o <= x"FFFFFFFF";
      when 3183 => data_o <= x"FFFFFFFF";
      when 3184 => data_o <= x"FFFFFFFF";
      when 3185 => data_o <= x"FFFFFFFF";
      when 3186 => data_o <= x"FFFFFFFF";
      when 3187 => data_o <= x"FFFFFFFF";
      when 3188 => data_o <= x"FFFFFFFF";
      when 3189 => data_o <= x"FFFFFFFF";
      when 3190 => data_o <= x"FFFFFFFF";
      when 3191 => data_o <= x"FFFFFFFF";
      when 3192 => data_o <= x"FFFFFFFF";
      when 3193 => data_o <= x"FFFFFFFF";
      when 3194 => data_o <= x"FFFFFFFF";
      when 3195 => data_o <= x"FFFFFFFF";
      when 3196 => data_o <= x"FFFFFFFF";
      when 3197 => data_o <= x"FFFFFFFF";
      when 3198 => data_o <= x"FFFFFFFF";
      when 3199 => data_o <= x"FFFFFFFF";
      when 3200 => data_o <= x"FFFFFFFF";
      when 3201 => data_o <= x"FFFFFFFF";
      when 3202 => data_o <= x"FFFFFFFF";
      when 3203 => data_o <= x"FFFFFFFF";
      when 3204 => data_o <= x"FFFFFFFF";
      when 3205 => data_o <= x"FFFFFFFF";
      when 3206 => data_o <= x"FFFFFFFF";
      when 3207 => data_o <= x"FFFFFFFF";
      when 3208 => data_o <= x"FFFFFFFF";
      when 3209 => data_o <= x"FFFFFFFF";
      when 3210 => data_o <= x"FFFFFFFF";
      when 3211 => data_o <= x"FFFFFFFF";
      when 3212 => data_o <= x"FFFFFFFF";
      when 3213 => data_o <= x"FFFFFFFF";
      when 3214 => data_o <= x"FFFFFFFF";
      when 3215 => data_o <= x"FFFFFFFF";
      when 3216 => data_o <= x"FFFFFFFF";
      when 3217 => data_o <= x"FFFFFFFF";
      when 3218 => data_o <= x"FFFFFFFF";
      when 3219 => data_o <= x"FFFFFFFF";
      when 3220 => data_o <= x"FFFFFFFF";
      when 3221 => data_o <= x"FFFFFFFF";
      when 3222 => data_o <= x"FFFFFFFF";
      when 3223 => data_o <= x"FFFFFFFF";
      when 3224 => data_o <= x"FFFFFFFF";
      when 3225 => data_o <= x"FFFFFFFF";
      when 3226 => data_o <= x"FFFFFFFF";
      when 3227 => data_o <= x"FFFFFFFF";
      when 3228 => data_o <= x"FFFFFFFF";
      when 3229 => data_o <= x"FFFFFFFF";
      when 3230 => data_o <= x"FFFFFFFF";
      when 3231 => data_o <= x"FFFFFFFF";
      when 3232 => data_o <= x"FFFFFFFF";
      when 3233 => data_o <= x"FFFFFFFF";
      when 3234 => data_o <= x"FFFFFFFF";
      when 3235 => data_o <= x"FFFFFFFF";
      when 3236 => data_o <= x"FFFFFFFF";
      when 3237 => data_o <= x"FFFFFFFF";
      when 3238 => data_o <= x"FFFFFFFF";
      when 3239 => data_o <= x"FFFFFFFF";
      when 3240 => data_o <= x"FFFFFFFF";
      when 3241 => data_o <= x"FFFFFFFF";
      when 3242 => data_o <= x"FFFFFFFF";
      when 3243 => data_o <= x"FFFFFFFF";
      when 3244 => data_o <= x"FFFFFFFF";
      when 3245 => data_o <= x"FFFFFFFF";
      when 3246 => data_o <= x"FFFFFFFF";
      when 3247 => data_o <= x"FFFFFFFF";
      when 3248 => data_o <= x"FFFFFFFF";
      when 3249 => data_o <= x"FFFFFFFF";
      when 3250 => data_o <= x"FFFFFFFF";
      when 3251 => data_o <= x"FFFFFFFF";
      when 3252 => data_o <= x"FFFFFFFF";
      when 3253 => data_o <= x"FFFFFFFF";
      when 3254 => data_o <= x"FFFFFFFF";
      when 3255 => data_o <= x"FFFFFFFF";
      when 3256 => data_o <= x"FFFFFFFF";
      when 3257 => data_o <= x"FFFFFFFF";
      when 3258 => data_o <= x"FFFFFFFF";
      when 3259 => data_o <= x"FFFFFFFF";
      when 3260 => data_o <= x"FFFFFFFF";
      when 3261 => data_o <= x"FFFFFFFF";
      when 3262 => data_o <= x"FFFFFFFF";
      when 3263 => data_o <= x"FFFFFFFF";
      when 3264 => data_o <= x"FFFFFFFF";
      when 3265 => data_o <= x"FFFFFFFF";
      when 3266 => data_o <= x"FFFFFFFF";
      when 3267 => data_o <= x"FFFFFFFF";
      when 3268 => data_o <= x"FFFFFFFF";
      when 3269 => data_o <= x"FFFFFFFF";
      when 3270 => data_o <= x"FFFFFFFF";
      when 3271 => data_o <= x"FFFFFFFF";
      when 3272 => data_o <= x"FFFFFFFF";
      when 3273 => data_o <= x"FFFFFFFF";
      when 3274 => data_o <= x"FFFFFFFF";
      when 3275 => data_o <= x"FFFFFFFF";
      when 3276 => data_o <= x"FFFFFFFF";
      when 3277 => data_o <= x"FFFFFFFF";
      when 3278 => data_o <= x"FFFFFFFF";
      when 3279 => data_o <= x"FFFFFFFF";
      when 3280 => data_o <= x"FFFFFFFF";
      when 3281 => data_o <= x"FFFFFFFF";
      when 3282 => data_o <= x"FFFFFFFF";
      when 3283 => data_o <= x"FFFFFFFF";
      when 3284 => data_o <= x"FFFFFFFF";
      when 3285 => data_o <= x"FFFFFFFF";
      when 3286 => data_o <= x"FFFFFFFF";
      when 3287 => data_o <= x"FFFFFFFF";
      when 3288 => data_o <= x"FFFFFFFF";
      when 3289 => data_o <= x"FFFFFFFF";
      when 3290 => data_o <= x"FFFFFFFF";
      when 3291 => data_o <= x"FFFFFFFF";
      when 3292 => data_o <= x"FFFFFFFF";
      when 3293 => data_o <= x"FFFFFFFF";
      when 3294 => data_o <= x"FFFFFFFF";
      when 3295 => data_o <= x"FFFFFFFF";
      when 3296 => data_o <= x"FFFFFFFF";
      when 3297 => data_o <= x"FFFFFFFF";
      when 3298 => data_o <= x"FFFFFFFF";
      when 3299 => data_o <= x"FFFFFFFF";
      when 3300 => data_o <= x"FFFFFFFF";
      when 3301 => data_o <= x"FFFFFFFF";
      when 3302 => data_o <= x"FFFFFFFF";
      when 3303 => data_o <= x"FFFFFFFF";
      when 3304 => data_o <= x"FFFFFFFF";
      when 3305 => data_o <= x"FFFFFFFF";
      when 3306 => data_o <= x"FFFFFFFF";
      when 3307 => data_o <= x"FFFFFFFF";
      when 3308 => data_o <= x"FFFFFFFF";
      when 3309 => data_o <= x"FFFFFFFF";
      when 3310 => data_o <= x"FFFFFFFF";
      when 3311 => data_o <= x"FFFFFFFF";
      when 3312 => data_o <= x"FFFFFFFF";
      when 3313 => data_o <= x"FFFFFFFF";
      when 3314 => data_o <= x"FFFFFFFF";
      when 3315 => data_o <= x"FFFFFFFF";
      when 3316 => data_o <= x"FFFFFFFF";
      when 3317 => data_o <= x"FFFFFFFF";
      when 3318 => data_o <= x"FFFFFFFF";
      when 3319 => data_o <= x"FFFFFFFF";
      when 3320 => data_o <= x"FFFFFFFF";
      when 3321 => data_o <= x"FFFFFFFF";
      when 3322 => data_o <= x"FFFFFFFF";
      when 3323 => data_o <= x"FFFFFFFF";
      when 3324 => data_o <= x"FFFFFFFF";
      when 3325 => data_o <= x"FFFFFFFF";
      when 3326 => data_o <= x"FFFFFFFF";
      when 3327 => data_o <= x"FFFFFFFF";
      when 3328 => data_o <= x"FFFFFFFF";
      when 3329 => data_o <= x"FFFFFFFF";
      when 3330 => data_o <= x"FFFFFFFF";
      when 3331 => data_o <= x"FFFFFFFF";
      when 3332 => data_o <= x"FFFFFFFF";
      when 3333 => data_o <= x"FFFFFFFF";
      when 3334 => data_o <= x"FFFFFFFF";
      when 3335 => data_o <= x"FFFFFFFF";
      when 3336 => data_o <= x"FFFFFFFF";
      when 3337 => data_o <= x"FFFFFFFF";
      when 3338 => data_o <= x"FFFFFFFF";
      when 3339 => data_o <= x"FFFFFFFF";
      when 3340 => data_o <= x"FFFFFFFF";
      when 3341 => data_o <= x"FFFFFFFF";
      when 3342 => data_o <= x"FFFFFFFF";
      when 3343 => data_o <= x"FFFFFFFF";
      when 3344 => data_o <= x"FFFFFFFF";
      when 3345 => data_o <= x"FFFFFFFF";
      when 3346 => data_o <= x"FFFFFFFF";
      when 3347 => data_o <= x"FFFFFFFF";
      when 3348 => data_o <= x"FFFFFFFF";
      when 3349 => data_o <= x"FFFFFFFF";
      when 3350 => data_o <= x"FFFFFFFF";
      when 3351 => data_o <= x"FFFFFFFF";
      when 3352 => data_o <= x"FFFFFFFF";
      when 3353 => data_o <= x"FFFFFFFF";
      when 3354 => data_o <= x"FFFFFFFF";
      when 3355 => data_o <= x"FFFFFFFF";
      when 3356 => data_o <= x"FFFFFFFF";
      when 3357 => data_o <= x"FFFFFFFF";
      when 3358 => data_o <= x"FFFFFFFF";
      when 3359 => data_o <= x"FFFFFFFF";
      when 3360 => data_o <= x"FFFFFFFF";
      when 3361 => data_o <= x"FFFFFFFF";
      when 3362 => data_o <= x"FFFFFFFF";
      when 3363 => data_o <= x"FFFFFFFF";
      when 3364 => data_o <= x"FFFFFFFF";
      when 3365 => data_o <= x"FFFFFFFF";
      when 3366 => data_o <= x"FFFFFFFF";
      when 3367 => data_o <= x"FFFFFFFF";
      when 3368 => data_o <= x"FFFFFFFF";
      when 3369 => data_o <= x"FFFFFFFF";
      when 3370 => data_o <= x"FFFFFFFF";
      when 3371 => data_o <= x"FFFFFFFF";
      when 3372 => data_o <= x"FFFFFFFF";
      when 3373 => data_o <= x"FFFFFFFF";
      when 3374 => data_o <= x"FFFFFFFF";
      when 3375 => data_o <= x"FFFFFFFF";
      when 3376 => data_o <= x"FFFFFFFF";
      when 3377 => data_o <= x"FFFFFFFF";
      when 3378 => data_o <= x"FFFFFFFF";
      when 3379 => data_o <= x"FFFFFFFF";
      when 3380 => data_o <= x"FFFFFFFF";
      when 3381 => data_o <= x"FFFFFFFF";
      when 3382 => data_o <= x"FFFFFFFF";
      when 3383 => data_o <= x"FFFFFFFF";
      when 3384 => data_o <= x"FFFFFFFF";
      when 3385 => data_o <= x"FFFFFFFF";
      when 3386 => data_o <= x"FFFFFFFF";
      when 3387 => data_o <= x"FFFFFFFF";
      when 3388 => data_o <= x"FFFFFFFF";
      when 3389 => data_o <= x"FFFFFFFF";
      when 3390 => data_o <= x"FFFFFFFF";
      when 3391 => data_o <= x"FFFFFFFF";
      when 3392 => data_o <= x"FFFFFFFF";
      when 3393 => data_o <= x"FFFFFFFF";
      when 3394 => data_o <= x"FFFFFFFF";
      when 3395 => data_o <= x"FFFFFFFF";
      when 3396 => data_o <= x"FFFFFFFF";
      when 3397 => data_o <= x"FFFFFFFF";
      when 3398 => data_o <= x"FFFFFFFF";
      when 3399 => data_o <= x"FFFFFFFF";
      when 3400 => data_o <= x"FFFFFFFF";
      when 3401 => data_o <= x"FFFFFFFF";
      when 3402 => data_o <= x"FFFFFFFF";
      when 3403 => data_o <= x"FFFFFFFF";
      when 3404 => data_o <= x"FFFFFFFF";
      when 3405 => data_o <= x"FFFFFFFF";
      when 3406 => data_o <= x"FFFFFFFF";
      when 3407 => data_o <= x"FFFFFFFF";
      when 3408 => data_o <= x"FFFFFFFF";
      when 3409 => data_o <= x"FFFFFFFF";
      when 3410 => data_o <= x"FFFFFFFF";
      when 3411 => data_o <= x"FFFFFFFF";
      when 3412 => data_o <= x"FFFFFFFF";
      when 3413 => data_o <= x"FFFFFFFF";
      when 3414 => data_o <= x"FFFFFFFF";
      when 3415 => data_o <= x"FFFFFFFF";
      when 3416 => data_o <= x"FFFFFFFF";
      when 3417 => data_o <= x"FFFFFFFF";
      when 3418 => data_o <= x"FFFFFFFF";
      when 3419 => data_o <= x"FFFFFFFF";
      when 3420 => data_o <= x"FFFFFFFF";
      when 3421 => data_o <= x"FFFFFFFF";
      when 3422 => data_o <= x"FFFFFFFF";
      when 3423 => data_o <= x"FFFFFFFF";
      when 3424 => data_o <= x"FFFFFFFF";
      when 3425 => data_o <= x"FFFFFFFF";
      when 3426 => data_o <= x"FFFFFFFF";
      when 3427 => data_o <= x"FFFFFFFF";
      when 3428 => data_o <= x"FFFFFFFF";
      when 3429 => data_o <= x"FFFFFFFF";
      when 3430 => data_o <= x"FFFFFFFF";
      when 3431 => data_o <= x"FFFFFFFF";
      when 3432 => data_o <= x"FFFFFFFF";
      when 3433 => data_o <= x"FFFFFFFF";
      when 3434 => data_o <= x"FFFFFFFF";
      when 3435 => data_o <= x"FFFFFFFF";
      when 3436 => data_o <= x"FFFFFFFF";
      when 3437 => data_o <= x"FFFFFFFF";
      when 3438 => data_o <= x"FFFFFFFF";
      when 3439 => data_o <= x"FFFFFFFF";
      when 3440 => data_o <= x"FFFFFFFF";
      when 3441 => data_o <= x"FFFFFFFF";
      when 3442 => data_o <= x"FFFFFFFF";
      when 3443 => data_o <= x"FFFFFFFF";
      when 3444 => data_o <= x"FFFFFFFF";
      when 3445 => data_o <= x"FFFFFFFF";
      when 3446 => data_o <= x"FFFFFFFF";
      when 3447 => data_o <= x"FFFFFFFF";
      when 3448 => data_o <= x"FFFFFFFF";
      when 3449 => data_o <= x"FFFFFFFF";
      when 3450 => data_o <= x"FFFFFFFF";
      when 3451 => data_o <= x"FFFFFFFF";
      when 3452 => data_o <= x"FFFFFFFF";
      when 3453 => data_o <= x"FFFFFFFF";
      when 3454 => data_o <= x"FFFFFFFF";
      when 3455 => data_o <= x"FFFFFFFF";
      when 3456 => data_o <= x"FFFFFFFF";
      when 3457 => data_o <= x"FFFFFFFF";
      when 3458 => data_o <= x"FFFFFFFF";
      when 3459 => data_o <= x"FFFFFFFF";
      when 3460 => data_o <= x"FFFFFFFF";
      when 3461 => data_o <= x"FFFFFFFF";
      when 3462 => data_o <= x"FFFFFFFF";
      when 3463 => data_o <= x"FFFFFFFF";
      when 3464 => data_o <= x"FFFFFFFF";
      when 3465 => data_o <= x"FFFFFFFF";
      when 3466 => data_o <= x"FFFFFFFF";
      when 3467 => data_o <= x"FFFFFFFF";
      when 3468 => data_o <= x"FFFFFFFF";
      when 3469 => data_o <= x"FFFFFFFF";
      when 3470 => data_o <= x"FFFFFFFF";
      when 3471 => data_o <= x"FFFFFFFF";
      when 3472 => data_o <= x"FFFFFFFF";
      when 3473 => data_o <= x"FFFFFFFF";
      when 3474 => data_o <= x"FFFFFFFF";
      when 3475 => data_o <= x"FFFFFFFF";
      when 3476 => data_o <= x"FFFFFFFF";
      when 3477 => data_o <= x"FFFFFFFF";
      when 3478 => data_o <= x"FFFFFFFF";
      when 3479 => data_o <= x"FFFFFFFF";
      when 3480 => data_o <= x"FFFFFFFF";
      when 3481 => data_o <= x"FFFFFFFF";
      when 3482 => data_o <= x"FFFFFFFF";
      when 3483 => data_o <= x"FFFFFFFF";
      when 3484 => data_o <= x"FFFFFFFF";
      when 3485 => data_o <= x"FFFFFFFF";
      when 3486 => data_o <= x"FFFFFFFF";
      when 3487 => data_o <= x"FFFFFFFF";
      when 3488 => data_o <= x"FFFFFFFF";
      when 3489 => data_o <= x"FFFFFFFF";
      when 3490 => data_o <= x"FFFFFFFF";
      when 3491 => data_o <= x"FFFFFFFF";
      when 3492 => data_o <= x"FFFFFFFF";
      when 3493 => data_o <= x"FFFFFFFF";
      when 3494 => data_o <= x"FFFFFFFF";
      when 3495 => data_o <= x"FFFFFFFF";
      when 3496 => data_o <= x"FFFFFFFF";
      when 3497 => data_o <= x"FFFFFFFF";
      when 3498 => data_o <= x"FFFFFFFF";
      when 3499 => data_o <= x"FFFFFFFF";
      when 3500 => data_o <= x"FFFFFFFF";
      when 3501 => data_o <= x"FFFFFFFF";
      when 3502 => data_o <= x"FFFFFFFF";
      when 3503 => data_o <= x"FFFFFFFF";
      when 3504 => data_o <= x"FFFFFFFF";
      when 3505 => data_o <= x"FFFFFFFF";
      when 3506 => data_o <= x"FFFFFFFF";
      when 3507 => data_o <= x"FFFFFFFF";
      when 3508 => data_o <= x"FFFFFFFF";
      when 3509 => data_o <= x"FFFFFFFF";
      when 3510 => data_o <= x"FFFFFFFF";
      when 3511 => data_o <= x"FFFFFFFF";
      when 3512 => data_o <= x"FFFFFFFF";
      when 3513 => data_o <= x"FFFFFFFF";
      when 3514 => data_o <= x"FFFFFFFF";
      when 3515 => data_o <= x"FFFFFFFF";
      when 3516 => data_o <= x"FFFFFFFF";
      when 3517 => data_o <= x"FFFFFFFF";
      when 3518 => data_o <= x"FFFFFFFF";
      when 3519 => data_o <= x"FFFFFFFF";
      when 3520 => data_o <= x"FFFFFFFF";
      when 3521 => data_o <= x"FFFFFFFF";
      when 3522 => data_o <= x"FFFFFFFF";
      when 3523 => data_o <= x"FFFFFFFF";
      when 3524 => data_o <= x"FFFFFFFF";
      when 3525 => data_o <= x"FFFFFFFF";
      when 3526 => data_o <= x"FFFFFFFF";
      when 3527 => data_o <= x"FFFFFFFF";
      when 3528 => data_o <= x"FFFFFFFF";
      when 3529 => data_o <= x"FFFFFFFF";
      when 3530 => data_o <= x"FFFFFFFF";
      when 3531 => data_o <= x"FFFFFFFF";
      when 3532 => data_o <= x"FFFFFFFF";
      when 3533 => data_o <= x"FFFFFFFF";
      when 3534 => data_o <= x"FFFFFFFF";
      when 3535 => data_o <= x"FFFFFFFF";
      when 3536 => data_o <= x"FFFFFFFF";
      when 3537 => data_o <= x"FFFFFFFF";
      when 3538 => data_o <= x"FFFFFFFF";
      when 3539 => data_o <= x"FFFFFFFF";
      when 3540 => data_o <= x"FFFFFFFF";
      when 3541 => data_o <= x"FFFFFFFF";
      when 3542 => data_o <= x"FFFFFFFF";
      when 3543 => data_o <= x"FFFFFFFF";
      when 3544 => data_o <= x"FFFFFFFF";
      when 3545 => data_o <= x"FFFFFFFF";
      when 3546 => data_o <= x"FFFFFFFF";
      when 3547 => data_o <= x"FFFFFFFF";
      when 3548 => data_o <= x"FFFFFFFF";
      when 3549 => data_o <= x"FFFFFFFF";
      when 3550 => data_o <= x"FFFFFFFF";
      when 3551 => data_o <= x"FFFFFFFF";
      when 3552 => data_o <= x"FFFFFFFF";
      when 3553 => data_o <= x"FFFFFFFF";
      when 3554 => data_o <= x"FFFFFFFF";
      when 3555 => data_o <= x"FFFFFFFF";
      when 3556 => data_o <= x"FFFFFFFF";
      when 3557 => data_o <= x"FFFFFFFF";
      when 3558 => data_o <= x"FFFFFFFF";
      when 3559 => data_o <= x"FFFFFFFF";
      when 3560 => data_o <= x"FFFFFFFF";
      when 3561 => data_o <= x"FFFFFFFF";
      when 3562 => data_o <= x"FFFFFFFF";
      when 3563 => data_o <= x"FFFFFFFF";
      when 3564 => data_o <= x"FFFFFFFF";
      when 3565 => data_o <= x"FFFFFFFF";
      when 3566 => data_o <= x"FFFFFFFF";
      when 3567 => data_o <= x"FFFFFFFF";
      when 3568 => data_o <= x"FFFFFFFF";
      when 3569 => data_o <= x"FFFFFFFF";
      when 3570 => data_o <= x"FFFFFFFF";
      when 3571 => data_o <= x"FFFFFFFF";
      when 3572 => data_o <= x"FFFFFFFF";
      when 3573 => data_o <= x"FFFFFFFF";
      when 3574 => data_o <= x"FFFFFFFF";
      when 3575 => data_o <= x"FFFFFFFF";
      when 3576 => data_o <= x"FFFFFFFF";
      when 3577 => data_o <= x"FFFFFFFF";
      when 3578 => data_o <= x"FFFFFFFF";
      when 3579 => data_o <= x"FFFFFFFF";
      when 3580 => data_o <= x"FFFFFFFF";
      when 3581 => data_o <= x"FFFFFFFF";
      when 3582 => data_o <= x"FFFFFFFF";
      when 3583 => data_o <= x"FFFFFFFF";
      when 3584 => data_o <= x"FFFFFFFF";
      when 3585 => data_o <= x"FFFFFFFF";
      when 3586 => data_o <= x"FFFFFFFF";
      when 3587 => data_o <= x"FFFFFFFF";
      when 3588 => data_o <= x"FFFFFFFF";
      when 3589 => data_o <= x"FFFFFFFF";
      when 3590 => data_o <= x"FFFFFFFF";
      when 3591 => data_o <= x"FFFFFFFF";
      when 3592 => data_o <= x"FFFFFFFF";
      when 3593 => data_o <= x"FFFFFFFF";
      when 3594 => data_o <= x"FFFFFFFF";
      when 3595 => data_o <= x"FFFFFFFF";
      when 3596 => data_o <= x"FFFFFFFF";
      when 3597 => data_o <= x"FFFFFFFF";
      when 3598 => data_o <= x"FFFFFFFF";
      when 3599 => data_o <= x"FFFFFFFF";
      when 3600 => data_o <= x"FFFFFFFF";
      when 3601 => data_o <= x"FFFFFFFF";
      when 3602 => data_o <= x"FFFFFFFF";
      when 3603 => data_o <= x"FFFFFFFF";
      when 3604 => data_o <= x"FFFFFFFF";
      when 3605 => data_o <= x"FFFFFFFF";
      when 3606 => data_o <= x"FFFFFFFF";
      when 3607 => data_o <= x"FFFFFFFF";
      when 3608 => data_o <= x"FFFFFFFF";
      when 3609 => data_o <= x"FFFFFFFF";
      when 3610 => data_o <= x"FFFFFFFF";
      when 3611 => data_o <= x"FFFFFFFF";
      when 3612 => data_o <= x"FFFFFFFF";
      when 3613 => data_o <= x"FFFFFFFF";
      when 3614 => data_o <= x"FFFFFFFF";
      when 3615 => data_o <= x"FFFFFFFF";
      when 3616 => data_o <= x"FFFFFFFF";
      when 3617 => data_o <= x"FFFFFFFF";
      when 3618 => data_o <= x"FFFFFFFF";
      when 3619 => data_o <= x"FFFFFFFF";
      when 3620 => data_o <= x"FFFFFFFF";
      when 3621 => data_o <= x"FFFFFFFF";
      when 3622 => data_o <= x"FFFFFFFF";
      when 3623 => data_o <= x"FFFFFFFF";
      when 3624 => data_o <= x"FFFFFFFF";
      when 3625 => data_o <= x"FFFFFFFF";
      when 3626 => data_o <= x"FFFFFFFF";
      when 3627 => data_o <= x"FFFFFFFF";
      when 3628 => data_o <= x"FFFFFFFF";
      when 3629 => data_o <= x"FFFFFFFF";
      when 3630 => data_o <= x"FFFFFFFF";
      when 3631 => data_o <= x"FFFFFFFF";
      when 3632 => data_o <= x"FFFFFFFF";
      when 3633 => data_o <= x"FFFFFFFF";
      when 3634 => data_o <= x"FFFFFFFF";
      when 3635 => data_o <= x"FFFFFFFF";
      when 3636 => data_o <= x"FFFFFFFF";
      when 3637 => data_o <= x"FFFFFFFF";
      when 3638 => data_o <= x"FFFFFFFF";
      when 3639 => data_o <= x"FFFFFFFF";
      when 3640 => data_o <= x"FFFFFFFF";
      when 3641 => data_o <= x"FFFFFFFF";
      when 3642 => data_o <= x"FFFFFFFF";
      when 3643 => data_o <= x"FFFFFFFF";
      when 3644 => data_o <= x"FFFFFFFF";
      when 3645 => data_o <= x"FFFFFFFF";
      when 3646 => data_o <= x"FFFFFFFF";
      when 3647 => data_o <= x"FFFFFFFF";
      when 3648 => data_o <= x"FFFFFFFF";
      when 3649 => data_o <= x"FFFFFFFF";
      when 3650 => data_o <= x"FFFFFFFF";
      when 3651 => data_o <= x"FFFFFFFF";
      when 3652 => data_o <= x"FFFFFFFF";
      when 3653 => data_o <= x"FFFFFFFF";
      when 3654 => data_o <= x"FFFFFFFF";
      when 3655 => data_o <= x"FFFFFFFF";
      when 3656 => data_o <= x"FFFFFFFF";
      when 3657 => data_o <= x"FFFFFFFF";
      when 3658 => data_o <= x"FFFFFFFF";
      when 3659 => data_o <= x"FFFFFFFF";
      when 3660 => data_o <= x"FFFFFFFF";
      when 3661 => data_o <= x"FFFFFFFF";
      when 3662 => data_o <= x"FFFFFFFF";
      when 3663 => data_o <= x"FFFFFFFF";
      when 3664 => data_o <= x"FFFFFFFF";
      when 3665 => data_o <= x"FFFFFFFF";
      when 3666 => data_o <= x"FFFFFFFF";
      when 3667 => data_o <= x"FFFFFFFF";
      when 3668 => data_o <= x"FFFFFFFF";
      when 3669 => data_o <= x"FFFFFFFF";
      when 3670 => data_o <= x"FFFFFFFF";
      when 3671 => data_o <= x"FFFFFFFF";
      when 3672 => data_o <= x"FFFFFFFF";
      when 3673 => data_o <= x"FFFFFFFF";
      when 3674 => data_o <= x"FFFFFFFF";
      when 3675 => data_o <= x"FFFFFFFF";
      when 3676 => data_o <= x"FFFFFFFF";
      when 3677 => data_o <= x"FFFFFFFF";
      when 3678 => data_o <= x"FFFFFFFF";
      when 3679 => data_o <= x"FFFFFFFF";
      when 3680 => data_o <= x"FFFFFFFF";
      when 3681 => data_o <= x"FFFFFFFF";
      when 3682 => data_o <= x"FFFFFFFF";
      when 3683 => data_o <= x"FFFFFFFF";
      when 3684 => data_o <= x"FFFFFFFF";
      when 3685 => data_o <= x"FFFFFFFF";
      when 3686 => data_o <= x"FFFFFFFF";
      when 3687 => data_o <= x"FFFFFFFF";
      when 3688 => data_o <= x"FFFFFFFF";
      when 3689 => data_o <= x"FFFFFFFF";
      when 3690 => data_o <= x"FFFFFFFF";
      when 3691 => data_o <= x"FFFFFFFF";
      when 3692 => data_o <= x"FFFFFFFF";
      when 3693 => data_o <= x"FFFFFFFF";
      when 3694 => data_o <= x"FFFFFFFF";
      when 3695 => data_o <= x"FFFFFFFF";
      when 3696 => data_o <= x"FFFFFFFF";
      when 3697 => data_o <= x"FFFFFFFF";
      when 3698 => data_o <= x"FFFFFFFF";
      when 3699 => data_o <= x"FFFFFFFF";
      when 3700 => data_o <= x"FFFFFFFF";
      when 3701 => data_o <= x"FFFFFFFF";
      when 3702 => data_o <= x"FFFFFFFF";
      when 3703 => data_o <= x"FFFFFFFF";
      when 3704 => data_o <= x"FFFFFFFF";
      when 3705 => data_o <= x"FFFFFFFF";
      when 3706 => data_o <= x"FFFFFFFF";
      when 3707 => data_o <= x"FFFFFFFF";
      when 3708 => data_o <= x"FFFFFFFF";
      when 3709 => data_o <= x"FFFFFFFF";
      when 3710 => data_o <= x"FFFFFFFF";
      when 3711 => data_o <= x"FFFFFFFF";
      when 3712 => data_o <= x"FFFFFFFF";
      when 3713 => data_o <= x"FFFFFFFF";
      when 3714 => data_o <= x"FFFFFFFF";
      when 3715 => data_o <= x"FFFFFFFF";
      when 3716 => data_o <= x"FFFFFFFF";
      when 3717 => data_o <= x"FFFFFFFF";
      when 3718 => data_o <= x"FFFFFFFF";
      when 3719 => data_o <= x"FFFFFFFF";
      when 3720 => data_o <= x"FFFFFFFF";
      when 3721 => data_o <= x"FFFFFFFF";
      when 3722 => data_o <= x"FFFFFFFF";
      when 3723 => data_o <= x"FFFFFFFF";
      when 3724 => data_o <= x"FFFFFFFF";
      when 3725 => data_o <= x"FFFFFFFF";
      when 3726 => data_o <= x"FFFFFFFF";
      when 3727 => data_o <= x"FFFFFFFF";
      when 3728 => data_o <= x"FFFFFFFF";
      when 3729 => data_o <= x"FFFFFFFF";
      when 3730 => data_o <= x"FFFFFFFF";
      when 3731 => data_o <= x"FFFFFFFF";
      when 3732 => data_o <= x"FFFFFFFF";
      when 3733 => data_o <= x"FFFFFFFF";
      when 3734 => data_o <= x"FFFFFFFF";
      when 3735 => data_o <= x"FFFFFFFF";
      when 3736 => data_o <= x"FFFFFFFF";
      when 3737 => data_o <= x"FFFFFFFF";
      when 3738 => data_o <= x"FFFFFFFF";
      when 3739 => data_o <= x"FFFFFFFF";
      when 3740 => data_o <= x"FFFFFFFF";
      when 3741 => data_o <= x"FFFFFFFF";
      when 3742 => data_o <= x"FFFFFFFF";
      when 3743 => data_o <= x"FFFFFFFF";
      when 3744 => data_o <= x"FFFFFFFF";
      when 3745 => data_o <= x"FFFFFFFF";
      when 3746 => data_o <= x"FFFFFFFF";
      when 3747 => data_o <= x"FFFFFFFF";
      when 3748 => data_o <= x"FFFFFFFF";
      when 3749 => data_o <= x"FFFFFFFF";
      when 3750 => data_o <= x"FFFFFFFF";
      when 3751 => data_o <= x"FFFFFFFF";
      when 3752 => data_o <= x"FFFFFFFF";
      when 3753 => data_o <= x"FFFFFFFF";
      when 3754 => data_o <= x"FFFFFFFF";
      when 3755 => data_o <= x"FFFFFFFF";
      when 3756 => data_o <= x"FFFFFFFF";
      when 3757 => data_o <= x"FFFFFFFF";
      when 3758 => data_o <= x"FFFFFFFF";
      when 3759 => data_o <= x"FFFFFFFF";
      when 3760 => data_o <= x"FFFFFFFF";
      when 3761 => data_o <= x"FFFFFFFF";
      when 3762 => data_o <= x"FFFFFFFF";
      when 3763 => data_o <= x"FFFFFFFF";
      when 3764 => data_o <= x"FFFFFFFF";
      when 3765 => data_o <= x"FFFFFFFF";
      when 3766 => data_o <= x"FFFFFFFF";
      when 3767 => data_o <= x"FFFFFFFF";
      when 3768 => data_o <= x"FFFFFFFF";
      when 3769 => data_o <= x"FFFFFFFF";
      when 3770 => data_o <= x"FFFFFFFF";
      when 3771 => data_o <= x"FFFFFFFF";
      when 3772 => data_o <= x"FFFFFFFF";
      when 3773 => data_o <= x"FFFFFFFF";
      when 3774 => data_o <= x"FFFFFFFF";
      when 3775 => data_o <= x"FFFFFFFF";
      when 3776 => data_o <= x"FFFFFFFF";
      when 3777 => data_o <= x"FFFFFFFF";
      when 3778 => data_o <= x"FFFFFFFF";
      when 3779 => data_o <= x"FFFFFFFF";
      when 3780 => data_o <= x"FFFFFFFF";
      when 3781 => data_o <= x"FFFFFFFF";
      when 3782 => data_o <= x"FFFFFFFF";
      when 3783 => data_o <= x"FFFFFFFF";
      when 3784 => data_o <= x"FFFFFFFF";
      when 3785 => data_o <= x"FFFFFFFF";
      when 3786 => data_o <= x"FFFFFFFF";
      when 3787 => data_o <= x"FFFFFFFF";
      when 3788 => data_o <= x"FFFFFFFF";
      when 3789 => data_o <= x"FFFFFFFF";
      when 3790 => data_o <= x"FFFFFFFF";
      when 3791 => data_o <= x"FFFFFFFF";
      when 3792 => data_o <= x"FFFFFFFF";
      when 3793 => data_o <= x"FFFFFFFF";
      when 3794 => data_o <= x"FFFFFFFF";
      when 3795 => data_o <= x"FFFFFFFF";
      when 3796 => data_o <= x"FFFFFFFF";
      when 3797 => data_o <= x"FFFFFFFF";
      when 3798 => data_o <= x"FFFFFFFF";
      when 3799 => data_o <= x"FFFFFFFF";
      when 3800 => data_o <= x"FFFFFFFF";
      when 3801 => data_o <= x"FFFFFFFF";
      when 3802 => data_o <= x"FFFFFFFF";
      when 3803 => data_o <= x"FFFFFFFF";
      when 3804 => data_o <= x"FFFFFFFF";
      when 3805 => data_o <= x"FFFFFFFF";
      when 3806 => data_o <= x"FFFFFFFF";
      when 3807 => data_o <= x"FFFFFFFF";
      when 3808 => data_o <= x"FFFFFFFF";
      when 3809 => data_o <= x"FFFFFFFF";
      when 3810 => data_o <= x"FFFFFFFF";
      when 3811 => data_o <= x"FFFFFFFF";
      when 3812 => data_o <= x"FFFFFFFF";
      when 3813 => data_o <= x"FFFFFFFF";
      when 3814 => data_o <= x"FFFFFFFF";
      when 3815 => data_o <= x"FFFFFFFF";
      when 3816 => data_o <= x"FFFFFFFF";
      when 3817 => data_o <= x"FFFFFFFF";
      when 3818 => data_o <= x"FFFFFFFF";
      when 3819 => data_o <= x"FFFFFFFF";
      when 3820 => data_o <= x"FFFFFFFF";
      when 3821 => data_o <= x"FFFFFFFF";
      when 3822 => data_o <= x"FFFFFFFF";
      when 3823 => data_o <= x"FFFFFFFF";
      when 3824 => data_o <= x"FFFFFFFF";
      when 3825 => data_o <= x"FFFFFFFF";
      when 3826 => data_o <= x"FFFFFFFF";
      when 3827 => data_o <= x"FFFFFFFF";
      when 3828 => data_o <= x"FFFFFFFF";
      when 3829 => data_o <= x"FFFFFFFF";
      when 3830 => data_o <= x"FFFFFFFF";
      when 3831 => data_o <= x"FFFFFFFF";
      when 3832 => data_o <= x"FFFFFFFF";
      when 3833 => data_o <= x"FFFFFFFF";
      when 3834 => data_o <= x"FFFFFFFF";
      when 3835 => data_o <= x"FFFFFFFF";
      when 3836 => data_o <= x"FFFFFFFF";
      when 3837 => data_o <= x"FFFFFFFF";
      when 3838 => data_o <= x"FFFFFFFF";
      when 3839 => data_o <= x"FFFFFFFF";
      when 3840 => data_o <= x"FFFFFFFF";
      when 3841 => data_o <= x"FFFFFFFF";
      when 3842 => data_o <= x"FFFFFFFF";
      when 3843 => data_o <= x"FFFFFFFF";
      when 3844 => data_o <= x"FFFFFFFF";
      when 3845 => data_o <= x"FFFFFFFF";
      when 3846 => data_o <= x"FFFFFFFF";
      when 3847 => data_o <= x"FFFFFFFF";
      when 3848 => data_o <= x"FFFFFFFF";
      when 3849 => data_o <= x"FFFFFFFF";
      when 3850 => data_o <= x"FFFFFFFF";
      when 3851 => data_o <= x"FFFFFFFF";
      when 3852 => data_o <= x"FFFFFFFF";
      when 3853 => data_o <= x"FFFFFFFF";
      when 3854 => data_o <= x"FFFFFFFF";
      when 3855 => data_o <= x"FFFFFFFF";
      when 3856 => data_o <= x"FFFFFFFF";
      when 3857 => data_o <= x"FFFFFFFF";
      when 3858 => data_o <= x"FFFFFFFF";
      when 3859 => data_o <= x"FFFFFFFF";
      when 3860 => data_o <= x"FFFFFFFF";
      when 3861 => data_o <= x"FFFFFFFF";
      when 3862 => data_o <= x"FFFFFFFF";
      when 3863 => data_o <= x"FFFFFFFF";
      when 3864 => data_o <= x"FFFFFFFF";
      when 3865 => data_o <= x"FFFFFFFF";
      when 3866 => data_o <= x"FFFFFFFF";
      when 3867 => data_o <= x"FFFFFFFF";
      when 3868 => data_o <= x"FFFFFFFF";
      when 3869 => data_o <= x"FFFFFFFF";
      when 3870 => data_o <= x"FFFFFFFF";
      when 3871 => data_o <= x"FFFFFFFF";
      when 3872 => data_o <= x"FFFFFFFF";
      when 3873 => data_o <= x"FFFFFFFF";
      when 3874 => data_o <= x"FFFFFFFF";
      when 3875 => data_o <= x"FFFFFFFF";
      when 3876 => data_o <= x"FFFFFFFF";
      when 3877 => data_o <= x"FFFFFFFF";
      when 3878 => data_o <= x"FFFFFFFF";
      when 3879 => data_o <= x"FFFFFFFF";
      when 3880 => data_o <= x"FFFFFFFF";
      when 3881 => data_o <= x"FFFFFFFF";
      when 3882 => data_o <= x"FFFFFFFF";
      when 3883 => data_o <= x"FFFFFFFF";
      when 3884 => data_o <= x"FFFFFFFF";
      when 3885 => data_o <= x"FFFFFFFF";
      when 3886 => data_o <= x"FFFFFFFF";
      when 3887 => data_o <= x"FFFFFFFF";
      when 3888 => data_o <= x"FFFFFFFF";
      when 3889 => data_o <= x"FFFFFFFF";
      when 3890 => data_o <= x"FFFFFFFF";
      when 3891 => data_o <= x"FFFFFFFF";
      when 3892 => data_o <= x"FFFFFFFF";
      when 3893 => data_o <= x"FFFFFFFF";
      when 3894 => data_o <= x"FFFFFFFF";
      when 3895 => data_o <= x"FFFFFFFF";
      when 3896 => data_o <= x"FFFFFFFF";
      when 3897 => data_o <= x"FFFFFFFF";
      when 3898 => data_o <= x"FFFFFFFF";
      when 3899 => data_o <= x"FFFFFFFF";
      when 3900 => data_o <= x"FFFFFFFF";
      when 3901 => data_o <= x"FFFFFFFF";
      when 3902 => data_o <= x"FFFFFFFF";
      when 3903 => data_o <= x"FFFFFFFF";
      when 3904 => data_o <= x"FFFFFFFF";
      when 3905 => data_o <= x"FFFFFFFF";
      when 3906 => data_o <= x"FFFFFFFF";
      when 3907 => data_o <= x"FFFFFFFF";
      when 3908 => data_o <= x"FFFFFFFF";
      when 3909 => data_o <= x"FFFFFFFF";
      when 3910 => data_o <= x"FFFFFFFF";
      when 3911 => data_o <= x"FFFFFFFF";
      when 3912 => data_o <= x"FFFFFFFF";
      when 3913 => data_o <= x"FFFFFFFF";
      when 3914 => data_o <= x"FFFFFFFF";
      when 3915 => data_o <= x"FFFFFFFF";
      when 3916 => data_o <= x"FFFFFFFF";
      when 3917 => data_o <= x"FFFFFFFF";
      when 3918 => data_o <= x"FFFFFFFF";
      when 3919 => data_o <= x"FFFFFFFF";
      when 3920 => data_o <= x"FFFFFFFF";
      when 3921 => data_o <= x"FFFFFFFF";
      when 3922 => data_o <= x"FFFFFFFF";
      when 3923 => data_o <= x"FFFFFFFF";
      when 3924 => data_o <= x"FFFFFFFF";
      when 3925 => data_o <= x"FFFFFFFF";
      when 3926 => data_o <= x"FFFFFFFF";
      when 3927 => data_o <= x"FFFFFFFF";
      when 3928 => data_o <= x"FFFFFFFF";
      when 3929 => data_o <= x"FFFFFFFF";
      when 3930 => data_o <= x"FFFFFFFF";
      when 3931 => data_o <= x"FFFFFFFF";
      when 3932 => data_o <= x"FFFFFFFF";
      when 3933 => data_o <= x"FFFFFFFF";
      when 3934 => data_o <= x"FFFFFFFF";
      when 3935 => data_o <= x"FFFFFFFF";
      when 3936 => data_o <= x"FFFFFFFF";
      when 3937 => data_o <= x"FFFFFFFF";
      when 3938 => data_o <= x"FFFFFFFF";
      when 3939 => data_o <= x"FFFFFFFF";
      when 3940 => data_o <= x"FFFFFFFF";
      when 3941 => data_o <= x"FFFFFFFF";
      when 3942 => data_o <= x"FFFFFFFF";
      when 3943 => data_o <= x"FFFFFFFF";
      when 3944 => data_o <= x"FFFFFFFF";
      when 3945 => data_o <= x"FFFFFFFF";
      when 3946 => data_o <= x"FFFFFFFF";
      when 3947 => data_o <= x"FFFFFFFF";
      when 3948 => data_o <= x"FFFFFFFF";
      when 3949 => data_o <= x"FFFFFFFF";
      when 3950 => data_o <= x"FFFFFFFF";
      when 3951 => data_o <= x"FFFFFFFF";
      when 3952 => data_o <= x"FFFFFFFF";
      when 3953 => data_o <= x"FFFFFFFF";
      when 3954 => data_o <= x"FFFFFFFF";
      when 3955 => data_o <= x"FFFFFFFF";
      when 3956 => data_o <= x"FFFFFFFF";
      when 3957 => data_o <= x"FFFFFFFF";
      when 3958 => data_o <= x"FFFFFFFF";
      when 3959 => data_o <= x"FFFFFFFF";
      when 3960 => data_o <= x"FFFFFFFF";
      when 3961 => data_o <= x"FFFFFFFF";
      when 3962 => data_o <= x"FFFFFFFF";
      when 3963 => data_o <= x"FFFFFFFF";
      when 3964 => data_o <= x"FFFFFFFF";
      when 3965 => data_o <= x"FFFFFFFF";
      when 3966 => data_o <= x"FFFFFFFF";
      when 3967 => data_o <= x"FFFFFFFF";
      when 3968 => data_o <= x"FFFFFFFF";
      when 3969 => data_o <= x"FFFFFFFF";
      when 3970 => data_o <= x"FFFFFFFF";
      when 3971 => data_o <= x"FFFFFFFF";
      when 3972 => data_o <= x"FFFFFFFF";
      when 3973 => data_o <= x"FFFFFFFF";
      when 3974 => data_o <= x"FFFFFFFF";
      when 3975 => data_o <= x"FFFFFFFF";
      when 3976 => data_o <= x"FFFFFFFF";
      when 3977 => data_o <= x"FFFFFFFF";
      when 3978 => data_o <= x"FFFFFFFF";
      when 3979 => data_o <= x"FFFFFFFF";
      when 3980 => data_o <= x"FFFFFFFF";
      when 3981 => data_o <= x"FFFFFFFF";
      when 3982 => data_o <= x"FFFFFFFF";
      when 3983 => data_o <= x"FFFFFFFF";
      when 3984 => data_o <= x"FFFFFFFF";
      when 3985 => data_o <= x"FFFFFFFF";
      when 3986 => data_o <= x"FFFFFFFF";
      when 3987 => data_o <= x"FFFFFFFF";
      when 3988 => data_o <= x"FFFFFFFF";
      when 3989 => data_o <= x"FFFFFFFF";
      when 3990 => data_o <= x"FFFFFFFF";
      when 3991 => data_o <= x"FFFFFFFF";
      when 3992 => data_o <= x"FFFFFFFF";
      when 3993 => data_o <= x"FFFFFFFF";
      when 3994 => data_o <= x"FFFFFFFF";
      when 3995 => data_o <= x"FFFFFFFF";
      when 3996 => data_o <= x"FFFFFFFF";
      when 3997 => data_o <= x"FFFFFFFF";
      when 3998 => data_o <= x"FFFFFFFF";
      when 3999 => data_o <= x"FFFFFFFF";
      when 4000 => data_o <= x"FFFFFFFF";
      when 4001 => data_o <= x"FFFFFFFF";
      when 4002 => data_o <= x"FFFFFFFF";
      when 4003 => data_o <= x"FFFFFFFF";
      when 4004 => data_o <= x"FFFFFFFF";
      when 4005 => data_o <= x"FFFFFFFF";
      when 4006 => data_o <= x"FFFFFFFF";
      when 4007 => data_o <= x"FFFFFFFF";
      when 4008 => data_o <= x"FFFFFFFF";
      when 4009 => data_o <= x"FFFFFFFF";
      when 4010 => data_o <= x"FFFFFFFF";
      when 4011 => data_o <= x"FFFFFFFF";
      when 4012 => data_o <= x"FFFFFFFF";
      when 4013 => data_o <= x"FFFFFFFF";
      when 4014 => data_o <= x"FFFFFFFF";
      when 4015 => data_o <= x"FFFFFFFF";
      when 4016 => data_o <= x"FFFFFFFF";
      when 4017 => data_o <= x"FFFFFFFF";
      when 4018 => data_o <= x"FFFFFFFF";
      when 4019 => data_o <= x"FFFFFFFF";
      when 4020 => data_o <= x"FFFFFFFF";
      when 4021 => data_o <= x"FFFFFFFF";
      when 4022 => data_o <= x"FFFFFFFF";
      when 4023 => data_o <= x"FFFFFFFF";
      when 4024 => data_o <= x"FFFFFFFF";
      when 4025 => data_o <= x"FFFFFFFF";
      when 4026 => data_o <= x"FFFFFFFF";
      when 4027 => data_o <= x"FFFFFFFF";
      when 4028 => data_o <= x"FFFFFFFF";
      when 4029 => data_o <= x"FFFFFFFF";
      when 4030 => data_o <= x"FFFFFFFF";
      when 4031 => data_o <= x"FFFFFFFF";
      when 4032 => data_o <= x"FFFFFFFF";
      when 4033 => data_o <= x"FFFFFFFF";
      when 4034 => data_o <= x"FFFFFFFF";
      when 4035 => data_o <= x"FFFFFFFF";
      when 4036 => data_o <= x"FFFFFFFF";
      when 4037 => data_o <= x"FFFFFFFF";
      when 4038 => data_o <= x"FFFFFFFF";
      when 4039 => data_o <= x"FFFFFFFF";
      when 4040 => data_o <= x"FFFFFFFF";
      when 4041 => data_o <= x"FFFFFFFF";
      when 4042 => data_o <= x"FFFFFFFF";
      when 4043 => data_o <= x"FFFFFFFF";
      when 4044 => data_o <= x"FFFFFFFF";
      when 4045 => data_o <= x"FFFFFFFF";
      when 4046 => data_o <= x"FFFFFFFF";
      when 4047 => data_o <= x"FFFFFFFF";
      when 4048 => data_o <= x"FFFFFFFF";
      when 4049 => data_o <= x"FFFFFFFF";
      when 4050 => data_o <= x"FFFFFFFF";
      when 4051 => data_o <= x"FFFFFFFF";
      when 4052 => data_o <= x"FFFFFFFF";
      when 4053 => data_o <= x"FFFFFFFF";
      when 4054 => data_o <= x"FFFFFFFF";
      when 4055 => data_o <= x"FFFFFFFF";
      when 4056 => data_o <= x"FFFFFFFF";
      when 4057 => data_o <= x"FFFFFFFF";
      when 4058 => data_o <= x"FFFFFFFF";
      when 4059 => data_o <= x"FFFFFFFF";
      when 4060 => data_o <= x"FFFFFFFF";
      when 4061 => data_o <= x"FFFFFFFF";
      when 4062 => data_o <= x"FFFFFFFF";
      when 4063 => data_o <= x"FFFFFFFF";
      when 4064 => data_o <= x"FFFFFFFF";
      when 4065 => data_o <= x"FFFFFFFF";
      when 4066 => data_o <= x"FFFFFFFF";
      when 4067 => data_o <= x"FFFFFFFF";
      when 4068 => data_o <= x"FFFFFFFF";
      when 4069 => data_o <= x"FFFFFFFF";
      when 4070 => data_o <= x"FFFFFFFF";
      when 4071 => data_o <= x"FFFFFFFF";
      when 4072 => data_o <= x"FFFFFFFF";
      when 4073 => data_o <= x"FFFFFFFF";
      when 4074 => data_o <= x"FFFFFFFF";
      when 4075 => data_o <= x"FFFFFFFF";
      when 4076 => data_o <= x"FFFFFFFF";
      when 4077 => data_o <= x"FFFFFFFF";
      when 4078 => data_o <= x"FFFFFFFF";
      when 4079 => data_o <= x"FFFFFFFF";
      when 4080 => data_o <= x"FFFFFFFF";
      when 4081 => data_o <= x"FFFFFFFF";
      when 4082 => data_o <= x"FFFFFFFF";
      when 4083 => data_o <= x"FFFFFFFF";
      when 4084 => data_o <= x"FFFFFFFF";
      when 4085 => data_o <= x"FFFFFFFF";
      when 4086 => data_o <= x"FFFFFFFF";
      when 4087 => data_o <= x"FFFFFFFF";
      when 4088 => data_o <= x"FFFFFFFF";
      when 4089 => data_o <= x"FFFFFFFF";
      when 4090 => data_o <= x"FFFFFFFF";
      when 4091 => data_o <= x"FFFFFFFF";
      when 4092 => data_o <= x"FFFFFFFF";
      when 4093 => data_o <= x"FFFFFFFF";
      when 4094 => data_o <= x"FFFFFFFF";
      when 4095 => data_o <= x"FFFFFFFF";
      when 4096 => data_o <= x"00004638";
      when 4097 => data_o <= x"12345678";
      when 4098 => data_o <= x"FEFFF334";
      when 4099 => data_o <= x"726F6605";
      when 4100 => data_o <= x"FFFF6874";
      when 4101 => data_o <= x"00FF0000";
      when 4102 => data_o <= x"0000146C";
      when 4103 => data_o <= x"000012E4";
      when 4104 => data_o <= x"FF000000";
      when 4105 => data_o <= x"FFFF7C01";
      when 4106 => data_o <= x"00000000";
      when 4107 => data_o <= x"00FF0000";
      when 4108 => data_o <= x"0000140C";
      when 4109 => data_o <= x"00001398";
      when 4110 => data_o <= x"FF004020";
      when 4111 => data_o <= x"706F6E03";
      when 4112 => data_o <= x"00000001";
      when 4113 => data_o <= x"00FF0000";
      when 4114 => data_o <= x"0000140C";
      when 4115 => data_o <= x"000012F4";
      when 4116 => data_o <= x"FF004038";
      when 4117 => data_o <= x"70756403";
      when 4118 => data_o <= x"00000003";
      when 4119 => data_o <= x"00FF0000";
      when 4120 => data_o <= x"0000140C";
      when 4121 => data_o <= x"000012F8";
      when 4122 => data_o <= x"FF004050";
      when 4123 => data_o <= x"FFFF2B01";
      when 4124 => data_o <= x"00000023";
      when 4125 => data_o <= x"00FF0000";
      when 4126 => data_o <= x"0000140C";
      when 4127 => data_o <= x"00001300";
      when 4128 => data_o <= x"FF004068";
      when 4129 => data_o <= x"FF2B6302";
      when 4130 => data_o <= x"00000012";
      when 4131 => data_o <= x"00FF0000";
      when 4132 => data_o <= x"0000140C";
      when 4133 => data_o <= x"00001304";
      when 4134 => data_o <= x"FF004080";
      when 4135 => data_o <= x"FF407202";
      when 4136 => data_o <= x"00000013";
      when 4137 => data_o <= x"00FF0000";
      when 4138 => data_o <= x"0000140C";
      when 4139 => data_o <= x"00001308";
      when 4140 => data_o <= x"FF004098";
      when 4141 => data_o <= x"646E6103";
      when 4142 => data_o <= x"00000039";
      when 4143 => data_o <= x"00FF0000";
      when 4144 => data_o <= x"0000140C";
      when 4145 => data_o <= x"0000130C";
      when 4146 => data_o <= x"FF0040B0";
      when 4147 => data_o <= x"65766F04";
      when 4148 => data_o <= x"FFFFFF72";
      when 4149 => data_o <= x"0000000A";
      when 4150 => data_o <= x"00FF0000";
      when 4151 => data_o <= x"0000140C";
      when 4152 => data_o <= x"00001310";
      when 4153 => data_o <= x"FF0040C8";
      when 4154 => data_o <= x"FF3E7202";
      when 4155 => data_o <= x"0000001B";
      when 4156 => data_o <= x"00FF0000";
      when 4157 => data_o <= x"0000140C";
      when 4158 => data_o <= x"00001314";
      when 4159 => data_o <= x"FF0040E4";
      when 4160 => data_o <= x"726F7803";
      when 4161 => data_o <= x"00000035";
      when 4162 => data_o <= x"00FF0000";
      when 4163 => data_o <= x"00001414";
      when 4164 => data_o <= x"000012E4";
      when 4165 => data_o <= x"FF0040FC";
      when 4166 => data_o <= x"73612103";
      when 4167 => data_o <= x"00000004";
      when 4168 => data_o <= x"00FF0000";
      when 4169 => data_o <= x"0000140C";
      when 4170 => data_o <= x"00001318";
      when 4171 => data_o <= x"FF004114";
      when 4172 => data_o <= x"FF2A3202";
      when 4173 => data_o <= x"0000000C";
      when 4174 => data_o <= x"00FF0000";
      when 4175 => data_o <= x"0000140C";
      when 4176 => data_o <= x"0000131C";
      when 4177 => data_o <= x"FF00412C";
      when 4178 => data_o <= x"632A3203";
      when 4179 => data_o <= x"0000000F";
      when 4180 => data_o <= x"00FF0000";
      when 4181 => data_o <= x"0000140C";
      when 4182 => data_o <= x"00001320";
      when 4183 => data_o <= x"FF004144";
      when 4184 => data_o <= x"2B216303";
      when 4185 => data_o <= x"0000000E";
      when 4186 => data_o <= x"00FF0000";
      when 4187 => data_o <= x"0000140C";
      when 4188 => data_o <= x"00001324";
      when 4189 => data_o <= x"FF00415C";
      when 4190 => data_o <= x"2B406303";
      when 4191 => data_o <= x"0000000E";
      when 4192 => data_o <= x"00FF0000";
      when 4193 => data_o <= x"0000140C";
      when 4194 => data_o <= x"00FFFFFD";
      when 4195 => data_o <= x"FF004174";
      when 4196 => data_o <= x"756F6305";
      when 4197 => data_o <= x"FFFF746E";
      when 4198 => data_o <= x"00000036";
      when 4199 => data_o <= x"00FF0000";
      when 4200 => data_o <= x"0000140C";
      when 4201 => data_o <= x"0000132C";
      when 4202 => data_o <= x"FF00418C";
      when 4203 => data_o <= x"FF406302";
      when 4204 => data_o <= x"00000017";
      when 4205 => data_o <= x"00FF0000";
      when 4206 => data_o <= x"0000140C";
      when 4207 => data_o <= x"00001330";
      when 4208 => data_o <= x"FF0041A8";
      when 4209 => data_o <= x"2B217703";
      when 4210 => data_o <= x"00000016";
      when 4211 => data_o <= x"00FF0000";
      when 4212 => data_o <= x"0000140C";
      when 4213 => data_o <= x"00001334";
      when 4214 => data_o <= x"FF0041C0";
      when 4215 => data_o <= x"2B407703";
      when 4216 => data_o <= x"0000001E";
      when 4217 => data_o <= x"00FF0000";
      when 4218 => data_o <= x"0000140C";
      when 4219 => data_o <= x"00001338";
      when 4220 => data_o <= x"FF0041D8";
      when 4221 => data_o <= x"FF407702";
      when 4222 => data_o <= x"00000027";
      when 4223 => data_o <= x"00FF0000";
      when 4224 => data_o <= x"0000140C";
      when 4225 => data_o <= x"0000133C";
      when 4226 => data_o <= x"FF0041F0";
      when 4227 => data_o <= x"FF2B2102";
      when 4228 => data_o <= x"00000026";
      when 4229 => data_o <= x"00FF0000";
      when 4230 => data_o <= x"0000140C";
      when 4231 => data_o <= x"00001340";
      when 4232 => data_o <= x"FF004208";
      when 4233 => data_o <= x"FF2B4002";
      when 4234 => data_o <= x"0000002E";
      when 4235 => data_o <= x"00FF0000";
      when 4236 => data_o <= x"0000140C";
      when 4237 => data_o <= x"00001344";
      when 4238 => data_o <= x"FF004220";
      when 4239 => data_o <= x"FFFF4001";
      when 4240 => data_o <= x"0000001C";
      when 4241 => data_o <= x"00FF0000";
      when 4242 => data_o <= x"0000140C";
      when 4243 => data_o <= x"00001348";
      when 4244 => data_o <= x"FF004238";
      when 4245 => data_o <= x"2F327503";
      when 4246 => data_o <= x"00000020";
      when 4247 => data_o <= x"00FF0000";
      when 4248 => data_o <= x"0000140C";
      when 4249 => data_o <= x"0000134C";
      when 4250 => data_o <= x"FF004250";
      when 4251 => data_o <= x"70657205";
      when 4252 => data_o <= x"FFFF6374";
      when 4253 => data_o <= x"00000028";
      when 4254 => data_o <= x"00FF0000";
      when 4255 => data_o <= x"0000140C";
      when 4256 => data_o <= x"00001350";
      when 4257 => data_o <= x"FF004268";
      when 4258 => data_o <= x"65722D05";
      when 4259 => data_o <= x"FFFF7470";
      when 4260 => data_o <= x"00000014";
      when 4261 => data_o <= x"00FF0000";
      when 4262 => data_o <= x"0000140C";
      when 4263 => data_o <= x"00001354";
      when 4264 => data_o <= x"FF004284";
      when 4265 => data_o <= x"FF2F3202";
      when 4266 => data_o <= x"00000019";
      when 4267 => data_o <= x"00FF0000";
      when 4268 => data_o <= x"0000140C";
      when 4269 => data_o <= x"00001358";
      when 4270 => data_o <= x"FF0042A0";
      when 4271 => data_o <= x"FF707302";
      when 4272 => data_o <= x"00000034";
      when 4273 => data_o <= x"00FF0000";
      when 4274 => data_o <= x"0000140C";
      when 4275 => data_o <= x"0000135C";
      when 4276 => data_o <= x"FF0042B8";
      when 4277 => data_o <= x"766E6906";
      when 4278 => data_o <= x"FF747265";
      when 4279 => data_o <= x"0000002F";
      when 4280 => data_o <= x"00FF0000";
      when 4281 => data_o <= x"0000140C";
      when 4282 => data_o <= x"00001360";
      when 4283 => data_o <= x"FF0042D0";
      when 4284 => data_o <= x"21707203";
      when 4285 => data_o <= x"00000011";
      when 4286 => data_o <= x"00FF0000";
      when 4287 => data_o <= x"0000140C";
      when 4288 => data_o <= x"00001364";
      when 4289 => data_o <= x"FF0042EC";
      when 4290 => data_o <= x"FF707202";
      when 4291 => data_o <= x"00000031";
      when 4292 => data_o <= x"00FF0000";
      when 4293 => data_o <= x"0000140C";
      when 4294 => data_o <= x"00001368";
      when 4295 => data_o <= x"FF004304";
      when 4296 => data_o <= x"726F7004";
      when 4297 => data_o <= x"FFFFFF74";
      when 4298 => data_o <= x"00000037";
      when 4299 => data_o <= x"00FF0000";
      when 4300 => data_o <= x"0000140C";
      when 4301 => data_o <= x"0000136C";
      when 4302 => data_o <= x"FF00431C";
      when 4303 => data_o <= x"21707303";
      when 4304 => data_o <= x"00000029";
      when 4305 => data_o <= x"00FF0000";
      when 4306 => data_o <= x"0000140C";
      when 4307 => data_o <= x"00001370";
      when 4308 => data_o <= x"FF004338";
      when 4309 => data_o <= x"FF707502";
      when 4310 => data_o <= x"0000003F";
      when 4311 => data_o <= x"00FF0000";
      when 4312 => data_o <= x"0000140C";
      when 4313 => data_o <= x"00001374";
      when 4314 => data_o <= x"FF004350";
      when 4315 => data_o <= x"21707503";
      when 4316 => data_o <= x"00000025";
      when 4317 => data_o <= x"00FF0000";
      when 4318 => data_o <= x"00001414";
      when 4319 => data_o <= x"000012E4";
      when 4320 => data_o <= x"FF004368";
      when 4321 => data_o <= x"74696C04";
      when 4322 => data_o <= x"FFFFFF78";
      when 4323 => data_o <= x"0000000D";
      when 4324 => data_o <= x"00FF0000";
      when 4325 => data_o <= x"00001414";
      when 4326 => data_o <= x"000012E4";
      when 4327 => data_o <= x"FF004380";
      when 4328 => data_o <= x"65737504";
      when 4329 => data_o <= x"FFFFFF72";
      when 4330 => data_o <= x"00000015";
      when 4331 => data_o <= x"00FF0000";
      when 4332 => data_o <= x"00001414";
      when 4333 => data_o <= x"000012E4";
      when 4334 => data_o <= x"FF00439C";
      when 4335 => data_o <= x"706D6A03";
      when 4336 => data_o <= x"0000002D";
      when 4337 => data_o <= x"00FF0000";
      when 4338 => data_o <= x"00001414";
      when 4339 => data_o <= x"000012E4";
      when 4340 => data_o <= x"FF0043B8";
      when 4341 => data_o <= x"73614003";
      when 4342 => data_o <= x"0000003D";
      when 4343 => data_o <= x"00FF0000";
      when 4344 => data_o <= x"00001414";
      when 4345 => data_o <= x"000012E4";
      when 4346 => data_o <= x"FF0043D0";
      when 4347 => data_o <= x"74696C03";
      when 4348 => data_o <= x"0000003B";
      when 4349 => data_o <= x"00FF0000";
      when 4350 => data_o <= x"0000140C";
      when 4351 => data_o <= x"00001378";
      when 4352 => data_o <= x"FF0043E8";
      when 4353 => data_o <= x"6F726404";
      when 4354 => data_o <= x"FFFFFF70";
      when 4355 => data_o <= x"0000001D";
      when 4356 => data_o <= x"00FF0000";
      when 4357 => data_o <= x"00001414";
      when 4358 => data_o <= x"000012E4";
      when 4359 => data_o <= x"FF004400";
      when 4360 => data_o <= x"6C616304";
      when 4361 => data_o <= x"FFFFFF6C";
      when 4362 => data_o <= x"00000009";
      when 4363 => data_o <= x"00FF0000";
      when 4364 => data_o <= x"0000140C";
      when 4365 => data_o <= x"0000137C";
      when 4366 => data_o <= x"FF00441C";
      when 4367 => data_o <= x"FF2B3102";
      when 4368 => data_o <= x"00000009";
      when 4369 => data_o <= x"00FF0000";
      when 4370 => data_o <= x"0000140C";
      when 4371 => data_o <= x"00001380";
      when 4372 => data_o <= x"FF004438";
      when 4373 => data_o <= x"61686305";
      when 4374 => data_o <= x"FFFF2B72";
      when 4375 => data_o <= x"00000021";
      when 4376 => data_o <= x"00FF0000";
      when 4377 => data_o <= x"0000140C";
      when 4378 => data_o <= x"00001384";
      when 4379 => data_o <= x"FF004450";
      when 4380 => data_o <= x"6C656305";
      when 4381 => data_o <= x"FFFF2B6C";
      when 4382 => data_o <= x"0000001F";
      when 4383 => data_o <= x"00FF0000";
      when 4384 => data_o <= x"0000140C";
      when 4385 => data_o <= x"00001388";
      when 4386 => data_o <= x"FF00446C";
      when 4387 => data_o <= x"FF723E02";
      when 4388 => data_o <= x"0000003C";
      when 4389 => data_o <= x"00FF0000";
      when 4390 => data_o <= x"0000140C";
      when 4391 => data_o <= x"0000138C";
      when 4392 => data_o <= x"FF004488";
      when 4393 => data_o <= x"61777304";
      when 4394 => data_o <= x"FFFFFF70";
      when 4395 => data_o <= x"00000008";
      when 4396 => data_o <= x"00FF0000";
      when 4397 => data_o <= x"00001440";
      when 4398 => data_o <= x"000012E4";
      when 4399 => data_o <= x"FF0044A0";
      when 4400 => data_o <= x"3A6F6E03";
      when 4401 => data_o <= x"00000038";
      when 4402 => data_o <= x"00FF0000";
      when 4403 => data_o <= x"00001440";
      when 4404 => data_o <= x"000012E4";
      when 4405 => data_o <= x"FF0044BC";
      when 4406 => data_o <= x"63666904";
      when 4407 => data_o <= x"FFFFFF3A";
      when 4408 => data_o <= x"0000003A";
      when 4409 => data_o <= x"00FF0000";
      when 4410 => data_o <= x"00001440";
      when 4411 => data_o <= x"000012E4";
      when 4412 => data_o <= x"FF0044D4";
      when 4413 => data_o <= x"7A666904";
      when 4414 => data_o <= x"FFFFFF3A";
      when 4415 => data_o <= x"00000030";
      when 4416 => data_o <= x"00FF0000";
      when 4417 => data_o <= x"00001440";
      when 4418 => data_o <= x"000012E4";
      when 4419 => data_o <= x"FF0044F0";
      when 4420 => data_o <= x"66692D04";
      when 4421 => data_o <= x"FFFFFF3A";
      when 4422 => data_o <= x"00000008";
      when 4423 => data_o <= x"00FF0000";
      when 4424 => data_o <= x"00001460";
      when 4425 => data_o <= x"000012E4";
      when 4426 => data_o <= x"FF00450C";
      when 4427 => data_o <= x"6F6E7C03";
      when 4428 => data_o <= x"00000038";
      when 4429 => data_o <= x"00FF0000";
      when 4430 => data_o <= x"00001460";
      when 4431 => data_o <= x"000012E4";
      when 4432 => data_o <= x"FF004528";
      when 4433 => data_o <= x"66697C04";
      when 4434 => data_o <= x"FFFFFF63";
      when 4435 => data_o <= x"0000003A";
      when 4436 => data_o <= x"00FF0000";
      when 4437 => data_o <= x"00001460";
      when 4438 => data_o <= x"000012E4";
      when 4439 => data_o <= x"FF004540";
      when 4440 => data_o <= x"66697C04";
      when 4441 => data_o <= x"FFFFFF7A";
      when 4442 => data_o <= x"00000030";
      when 4443 => data_o <= x"00FF0000";
      when 4444 => data_o <= x"00001460";
      when 4445 => data_o <= x"000012E4";
      when 4446 => data_o <= x"FF00455C";
      when 4447 => data_o <= x"692D7C04";
      when 4448 => data_o <= x"FFFFFF66";
      when 4449 => data_o <= x"00000024";
      when 4450 => data_o <= x"00FF0000";
      when 4451 => data_o <= x"0000140C";
      when 4452 => data_o <= x"00001390";
      when 4453 => data_o <= x"FF004578";
      when 4454 => data_o <= x"FF3D3002";
      when 4455 => data_o <= x"0000002C";
      when 4456 => data_o <= x"00FF0000";
      when 4457 => data_o <= x"0000140C";
      when 4458 => data_o <= x"00001394";
      when 4459 => data_o <= x"FF004594";
      when 4460 => data_o <= x"FF3C3002";
      when 4461 => data_o <= x"00000000";
      when 4462 => data_o <= x"00FF0000";
      when 4463 => data_o <= x"00001474";
      when 4464 => data_o <= x"000012EC";
      when 4465 => data_o <= x"FF0045AC";
      when 4466 => data_o <= x"61747306";
      when 4467 => data_o <= x"FF737574";
      when 4468 => data_o <= x"00000004";
      when 4469 => data_o <= x"00FF0000";
      when 4470 => data_o <= x"00001474";
      when 4471 => data_o <= x"000012EC";
      when 4472 => data_o <= x"FF0045C4";
      when 4473 => data_o <= x"6C6F6608";
      when 4474 => data_o <= x"65776F6C";
      when 4475 => data_o <= x"FFFFFF72";
      when 4476 => data_o <= x"00000008";
      when 4477 => data_o <= x"00FF0000";
      when 4478 => data_o <= x"00001474";
      when 4479 => data_o <= x"000012EC";
      when 4480 => data_o <= x"FF0045E0";
      when 4481 => data_o <= x"30707203";
      when 4482 => data_o <= x"0000000C";
      when 4483 => data_o <= x"00FF0000";
      when 4484 => data_o <= x"00001474";
      when 4485 => data_o <= x"000012EC";
      when 4486 => data_o <= x"FF004600";
      when 4487 => data_o <= x"30707303";
      when 4488 => data_o <= x"00000010";
      when 4489 => data_o <= x"00FF0000";
      when 4490 => data_o <= x"00001474";
      when 4491 => data_o <= x"000012EC";
      when 4492 => data_o <= x"FF004618";
      when 4493 => data_o <= x"736F7403";
      when 4494 => data_o <= x"000046D4";
      when 4495 => data_o <= x"69616D06";
      when 4496 => data_o <= x"FF662E6E";
      when 4497 => data_o <= x"00000004";
      when 4498 => data_o <= x"00FF0000";
      when 4499 => data_o <= x"070012BC";
      when 4500 => data_o <= x"000012B8";
      when 4501 => data_o <= x"FF004630";
      when 4502 => data_o <= x"6D75440B";
      when 4503 => data_o <= x"6C6F4370";
      when 4504 => data_o <= x"736E6D75";
      when 4505 => data_o <= x"00FF0001";
      when 4506 => data_o <= x"090012AC";
      when 4507 => data_o <= x"00000000";
      when 4508 => data_o <= x"FF004654";
      when 4509 => data_o <= x"6C6F63C8";
      when 4510 => data_o <= x"6F6F6264";
      when 4511 => data_o <= x"FFFFFF74";
      when 4512 => data_o <= x"00FF0001";
      when 4513 => data_o <= x"0A0012AC";
      when 4514 => data_o <= x"00000004";
      when 4515 => data_o <= x"FF004670";
      when 4516 => data_o <= x"666173C8";
      when 4517 => data_o <= x"646F6D65";
      when 4518 => data_o <= x"FFFFFF65";
      when 4519 => data_o <= x"00FF0001";
      when 4520 => data_o <= x"0B0012AC";
      when 4521 => data_o <= x"00000008";
      when 4522 => data_o <= x"FF00468C";
      when 4523 => data_o <= x"727265C8";
      when 4524 => data_o <= x"5349726F";
      when 4525 => data_o <= x"FFFFFF52";
      when 4526 => data_o <= x"00000001";
      when 4527 => data_o <= x"00FF0000";
      when 4528 => data_o <= x"0E0012BC";
      when 4529 => data_o <= x"000012B8";
      when 4530 => data_o <= x"FF0046A8";
      when 4531 => data_o <= x"74706F07";
      when 4532 => data_o <= x"736E6F69";
      when 4533 => data_o <= x"00004F00";
      when 4534 => data_o <= x"2F2E2E12";
      when 4535 => data_o <= x"662F2E2E";
      when 4536 => data_o <= x"6874726F";
      when 4537 => data_o <= x"726F632F";
      when 4538 => data_o <= x"FF662E65";
      when 4539 => data_o <= x"00000000";
      when 4540 => data_o <= x"01FF0000";
      when 4541 => data_o <= x"030012BC";
      when 4542 => data_o <= x"000012B8";
      when 4543 => data_o <= x"FF0046C8";
      when 4544 => data_o <= x"6C616605";
      when 4545 => data_o <= x"FFFF6573";
      when 4546 => data_o <= x"FFFFFFFF";
      when 4547 => data_o <= x"01FF0000";
      when 4548 => data_o <= x"040012BC";
      when 4549 => data_o <= x"000012B8";
      when 4550 => data_o <= x"FF0046FC";
      when 4551 => data_o <= x"75727404";
      when 4552 => data_o <= x"FFFFFF65";
      when 4553 => data_o <= x"00000020";
      when 4554 => data_o <= x"01FF0000";
      when 4555 => data_o <= x"050012BC";
      when 4556 => data_o <= x"000012B8";
      when 4557 => data_o <= x"FF004718";
      when 4558 => data_o <= x"FF6C6202";
      when 4559 => data_o <= x"01FF0001";
      when 4560 => data_o <= x"070012A8";
      when 4561 => data_o <= x"000012FC";
      when 4562 => data_o <= x"FF004734";
      when 4563 => data_o <= x"FFFF2DC1";
      when 4564 => data_o <= x"01FF0001";
      when 4565 => data_o <= x"080012A8";
      when 4566 => data_o <= x"00000018";
      when 4567 => data_o <= x"FF004748";
      when 4568 => data_o <= x"FFFF21C1";
      when 4569 => data_o <= x"01FF0001";
      when 4570 => data_o <= x"090012A8";
      when 4571 => data_o <= x"0000001C";
      when 4572 => data_o <= x"FF00475C";
      when 4573 => data_o <= x"FF2163C2";
      when 4574 => data_o <= x"01FF0001";
      when 4575 => data_o <= x"0A0012A8";
      when 4576 => data_o <= x"00000020";
      when 4577 => data_o <= x"FF004770";
      when 4578 => data_o <= x"FF2177C2";
      when 4579 => data_o <= x"01FF0002";
      when 4580 => data_o <= x"0B0012AC";
      when 4581 => data_o <= x"00000024";
      when 4582 => data_o <= x"FF004784";
      when 4583 => data_o <= x"FF212BC2";
      when 4584 => data_o <= x"01FF0002";
      when 4585 => data_o <= x"0C0012AC";
      when 4586 => data_o <= x"0000002C";
      when 4587 => data_o <= x"FF004798";
      when 4588 => data_o <= x"212B63C3";
      when 4589 => data_o <= x"01FF0001";
      when 4590 => data_o <= x"0D0012A8";
      when 4591 => data_o <= x"00000034";
      when 4592 => data_o <= x"FF0047AC";
      when 4593 => data_o <= x"67656EC6";
      when 4594 => data_o <= x"FF657461";
      when 4595 => data_o <= x"01FF0001";
      when 4596 => data_o <= x"0E0012A8";
      when 4597 => data_o <= x"00000038";
      when 4598 => data_o <= x"FF0047C0";
      when 4599 => data_o <= x"FF2D31C2";
      when 4600 => data_o <= x"01FF0001";
      when 4601 => data_o <= x"0F0012A8";
      when 4602 => data_o <= x"0000003C";
      when 4603 => data_o <= x"FF0047D8";
      when 4604 => data_o <= x"6C6563C5";
      when 4605 => data_o <= x"FFFF2D6C";
      when 4606 => data_o <= x"01FF0001";
      when 4607 => data_o <= x"100012A8";
      when 4608 => data_o <= x"00000040";
      when 4609 => data_o <= x"FF0047EC";
      when 4610 => data_o <= x"6C6563C5";
      when 4611 => data_o <= x"FFFF736C";
      when 4612 => data_o <= x"01FF0001";
      when 4613 => data_o <= x"110012A8";
      when 4614 => data_o <= x"00000044";
      when 4615 => data_o <= x"FF004804";
      when 4616 => data_o <= x"746F72C3";
      when 4617 => data_o <= x"01FF0001";
      when 4618 => data_o <= x"120012A8";
      when 4619 => data_o <= x"00000048";
      when 4620 => data_o <= x"FF00481C";
      when 4621 => data_o <= x"6F722DC4";
      when 4622 => data_o <= x"FFFFFF74";
      when 4623 => data_o <= x"01FF0001";
      when 4624 => data_o <= x"130012A8";
      when 4625 => data_o <= x"0000004C";
      when 4626 => data_o <= x"FF004830";
      when 4627 => data_o <= x"637574C4";
      when 4628 => data_o <= x"FFFFFF6B";
      when 4629 => data_o <= x"01FF0001";
      when 4630 => data_o <= x"140012A8";
      when 4631 => data_o <= x"00000050";
      when 4632 => data_o <= x"FF004848";
      when 4633 => data_o <= x"70696EC3";
      when 4634 => data_o <= x"01FF0002";
      when 4635 => data_o <= x"150012AC";
      when 4636 => data_o <= x"00000054";
      when 4637 => data_o <= x"FF004860";
      when 4638 => data_o <= x"723E3243";
      when 4639 => data_o <= x"01FF0002";
      when 4640 => data_o <= x"170012AC";
      when 4641 => data_o <= x"0000005C";
      when 4642 => data_o <= x"FF004874";
      when 4643 => data_o <= x"3E723243";
      when 4644 => data_o <= x"01FF0002";
      when 4645 => data_o <= x"190012AC";
      when 4646 => data_o <= x"00000064";
      when 4647 => data_o <= x"FF004888";
      when 4648 => data_o <= x"40723243";
      when 4649 => data_o <= x"01FF0001";
      when 4650 => data_o <= x"1B0012A8";
      when 4651 => data_o <= x"0000006C";
      when 4652 => data_o <= x"FF00489C";
      when 4653 => data_o <= x"726432C5";
      when 4654 => data_o <= x"FFFF706F";
      when 4655 => data_o <= x"01FF0001";
      when 4656 => data_o <= x"1C0012A8";
      when 4657 => data_o <= x"00000070";
      when 4658 => data_o <= x"FF0048B0";
      when 4659 => data_o <= x"756432C4";
      when 4660 => data_o <= x"FFFFFF70";
      when 4661 => data_o <= x"01FF0002";
      when 4662 => data_o <= x"1D0012AC";
      when 4663 => data_o <= x"00000074";
      when 4664 => data_o <= x"FF0048C8";
      when 4665 => data_o <= x"777332C5";
      when 4666 => data_o <= x"FFFF7061";
      when 4667 => data_o <= x"01FF0002";
      when 4668 => data_o <= x"1E0012AC";
      when 4669 => data_o <= x"0000007C";
      when 4670 => data_o <= x"FF0048E0";
      when 4671 => data_o <= x"766F32C5";
      when 4672 => data_o <= x"FFFF7265";
      when 4673 => data_o <= x"01FF0001";
      when 4674 => data_o <= x"1F0012A8";
      when 4675 => data_o <= x"00000084";
      when 4676 => data_o <= x"FF0048F8";
      when 4677 => data_o <= x"726433C5";
      when 4678 => data_o <= x"FFFF706F";
      when 4679 => data_o <= x"01FF0002";
      when 4680 => data_o <= x"200012AC";
      when 4681 => data_o <= x"00000088";
      when 4682 => data_o <= x"FF004910";
      when 4683 => data_o <= x"75643FC4";
      when 4684 => data_o <= x"FFFFFF70";
      when 4685 => data_o <= x"01FF0002";
      when 4686 => data_o <= x"210012AC";
      when 4687 => data_o <= x"00000090";
      when 4688 => data_o <= x"FF004928";
      when 4689 => data_o <= x"643E73C3";
      when 4690 => data_o <= x"01FF0001";
      when 4691 => data_o <= x"230012A8";
      when 4692 => data_o <= x"00000098";
      when 4693 => data_o <= x"FF004940";
      when 4694 => data_o <= x"746F6EC3";
      when 4695 => data_o <= x"01FF0001";
      when 4696 => data_o <= x"240012A8";
      when 4697 => data_o <= x"0000009C";
      when 4698 => data_o <= x"FF004954";
      when 4699 => data_o <= x"FFFF3DC1";
      when 4700 => data_o <= x"01FF0001";
      when 4701 => data_o <= x"250012A8";
      when 4702 => data_o <= x"000000A0";
      when 4703 => data_o <= x"FF004968";
      when 4704 => data_o <= x"FF3E3CC2";
      when 4705 => data_o <= x"01FF0001";
      when 4706 => data_o <= x"260012A8";
      when 4707 => data_o <= x"000000A4";
      when 4708 => data_o <= x"FF00497C";
      when 4709 => data_o <= x"3E3C30C3";
      when 4710 => data_o <= x"01FF0001";
      when 4711 => data_o <= x"270012A8";
      when 4712 => data_o <= x"000000A8";
      when 4713 => data_o <= x"FF004990";
      when 4714 => data_o <= x"FF3E30C2";
      when 4715 => data_o <= x"01FF0002";
      when 4716 => data_o <= x"280012AC";
      when 4717 => data_o <= x"000000AC";
      when 4718 => data_o <= x"FF0049A4";
      when 4719 => data_o <= x"696C61C7";
      when 4720 => data_o <= x"64656E67";
      when 4721 => data_o <= x"01FF0001";
      when 4722 => data_o <= x"290012AC";
      when 4723 => data_o <= x"000000B4";
      when 4724 => data_o <= x"FF0049B8";
      when 4725 => data_o <= x"FF4032C2";
      when 4726 => data_o <= x"01FF0001";
      when 4727 => data_o <= x"2A0012A8";
      when 4728 => data_o <= x"000000B8";
      when 4729 => data_o <= x"FF0049D0";
      when 4730 => data_o <= x"FF2132C2";
      when 4731 => data_o <= x"01FF0002";
      when 4732 => data_o <= x"2B0012AC";
      when 4733 => data_o <= x"000000BC";
      when 4734 => data_o <= x"FF0049E4";
      when 4735 => data_o <= x"736261C3";
      when 4736 => data_o <= x"01FF0001";
      when 4737 => data_o <= x"2C0012AC";
      when 4738 => data_o <= x"000000C4";
      when 4739 => data_o <= x"FF0049F8";
      when 4740 => data_o <= x"FF726FC2";
      when 4741 => data_o <= x"01FF0001";
      when 4742 => data_o <= x"2D0012AC";
      when 4743 => data_o <= x"000000C8";
      when 4744 => data_o <= x"FF004A0C";
      when 4745 => data_o <= x"657865C7";
      when 4746 => data_o <= x"65747563";
      when 4747 => data_o <= x"01FF0002";
      when 4748 => data_o <= x"2E0012AC";
      when 4749 => data_o <= x"000000CC";
      when 4750 => data_o <= x"FF004A20";
      when 4751 => data_o <= x"FF2B64C2";
      when 4752 => data_o <= x"01FF0003";
      when 4753 => data_o <= x"2F0012AC";
      when 4754 => data_o <= x"000000D4";
      when 4755 => data_o <= x"FF004A38";
      when 4756 => data_o <= x"656E64C7";
      when 4757 => data_o <= x"65746167";
      when 4758 => data_o <= x"01FF0002";
      when 4759 => data_o <= x"340012AC";
      when 4760 => data_o <= x"000000E0";
      when 4761 => data_o <= x"FF004A4C";
      when 4762 => data_o <= x"626164C4";
      when 4763 => data_o <= x"FFFFFF73";
      when 4764 => data_o <= x"01FF0001";
      when 4765 => data_o <= x"350012A8";
      when 4766 => data_o <= x"00001328";
      when 4767 => data_o <= x"FF004A64";
      when 4768 => data_o <= x"756F63C5";
      when 4769 => data_o <= x"FFFF746E";
      when 4770 => data_o <= x"01FF0002";
      when 4771 => data_o <= x"360012AC";
      when 4772 => data_o <= x"000000EC";
      when 4773 => data_o <= x"FF004A7C";
      when 4774 => data_o <= x"696874C5";
      when 4775 => data_o <= x"FFFF6472";
      when 4776 => data_o <= x"01FF0002";
      when 4777 => data_o <= x"370012AC";
      when 4778 => data_o <= x"000000F4";
      when 4779 => data_o <= x"FF004A94";
      when 4780 => data_o <= x"756F66C6";
      when 4781 => data_o <= x"FF687472";
      when 4782 => data_o <= x"01FF0004";
      when 4783 => data_o <= x"380012AC";
      when 4784 => data_o <= x"000000FC";
      when 4785 => data_o <= x"FF004AAC";
      when 4786 => data_o <= x"706564C5";
      when 4787 => data_o <= x"FFFF6874";
      when 4788 => data_o <= x"01FF0002";
      when 4789 => data_o <= x"390012AC";
      when 4790 => data_o <= x"0000010C";
      when 4791 => data_o <= x"FF004AC4";
      when 4792 => data_o <= x"636970C4";
      when 4793 => data_o <= x"FFFFFF6B";
      when 4794 => data_o <= x"01FF0003";
      when 4795 => data_o <= x"3A0012AC";
      when 4796 => data_o <= x"00000114";
      when 4797 => data_o <= x"FF004ADC";
      when 4798 => data_o <= x"636564C7";
      when 4799 => data_o <= x"6C616D69";
      when 4800 => data_o <= x"01FF0003";
      when 4801 => data_o <= x"3B0012AC";
      when 4802 => data_o <= x"00000120";
      when 4803 => data_o <= x"FF004AF4";
      when 4804 => data_o <= x"786568C3";
      when 4805 => data_o <= x"01FF0003";
      when 4806 => data_o <= x"3C0012AC";
      when 4807 => data_o <= x"0000012C";
      when 4808 => data_o <= x"FF004B0C";
      when 4809 => data_o <= x"6E696CC5";
      when 4810 => data_o <= x"FFFF3E6B";
      when 4811 => data_o <= x"01FF0005";
      when 4812 => data_o <= x"3F0012AC";
      when 4813 => data_o <= x"00000138";
      when 4814 => data_o <= x"FF004B20";
      when 4815 => data_o <= x"643F2845";
      when 4816 => data_o <= x"FFFF296F";
      when 4817 => data_o <= x"01FF0004";
      when 4818 => data_o <= x"440012AC";
      when 4819 => data_o <= x"0000014C";
      when 4820 => data_o <= x"FF004B38";
      when 4821 => data_o <= x"6F6C2846";
      when 4822 => data_o <= x"FF29706F";
      when 4823 => data_o <= x"01FF0006";
      when 4824 => data_o <= x"490012AC";
      when 4825 => data_o <= x"0000015C";
      when 4826 => data_o <= x"FF004B50";
      when 4827 => data_o <= x"6C2B2847";
      when 4828 => data_o <= x"29706F6F";
      when 4829 => data_o <= x"01FF0002";
      when 4830 => data_o <= x"510012AC";
      when 4831 => data_o <= x"00000174";
      when 4832 => data_o <= x"FF004B68";
      when 4833 => data_o <= x"FFFF6A41";
      when 4834 => data_o <= x"01FF0002";
      when 4835 => data_o <= x"520012AC";
      when 4836 => data_o <= x"0000017C";
      when 4837 => data_o <= x"FF004B80";
      when 4838 => data_o <= x"6C6E7546";
      when 4839 => data_o <= x"FF706F6F";
      when 4840 => data_o <= x"01FF0003";
      when 4841 => data_o <= x"550012AC";
      when 4842 => data_o <= x"00000184";
      when 4843 => data_o <= x"FF004B94";
      when 4844 => data_o <= x"666F2844";
      when 4845 => data_o <= x"FFFFFF29";
      when 4846 => data_o <= x"01FF0003";
      when 4847 => data_o <= x"5A0012AC";
      when 4848 => data_o <= x"00000190";
      when 4849 => data_o <= x"FF004BAC";
      when 4850 => data_o <= x"6F662845";
      when 4851 => data_o <= x"FFFF2972";
      when 4852 => data_o <= x"01FF0003";
      when 4853 => data_o <= x"600012AC";
      when 4854 => data_o <= x"0000019C";
      when 4855 => data_o <= x"FF004BC4";
      when 4856 => data_o <= x"74732848";
      when 4857 => data_o <= x"676E6972";
      when 4858 => data_o <= x"FFFFFF29";
      when 4859 => data_o <= x"01FF0002";
      when 4860 => data_o <= x"660012AC";
      when 4861 => data_o <= x"000001A8";
      when 4862 => data_o <= x"FF004BDC";
      when 4863 => data_o <= x"FF3C75C2";
      when 4864 => data_o <= x"01FF0001";
      when 4865 => data_o <= x"670012AC";
      when 4866 => data_o <= x"000001B0";
      when 4867 => data_o <= x"FF004BF8";
      when 4868 => data_o <= x"FF3E75C2";
      when 4869 => data_o <= x"01FF0003";
      when 4870 => data_o <= x"730012AC";
      when 4871 => data_o <= x"000001B4";
      when 4872 => data_o <= x"FF004C0C";
      when 4873 => data_o <= x"FFFF3CC1";
      when 4874 => data_o <= x"01FF0001";
      when 4875 => data_o <= x"780012AC";
      when 4876 => data_o <= x"000001C0";
      when 4877 => data_o <= x"FF004C20";
      when 4878 => data_o <= x"FFFF3EC1";
      when 4879 => data_o <= x"01FF0006";
      when 4880 => data_o <= x"7A0012AC";
      when 4881 => data_o <= x"000001C4";
      when 4882 => data_o <= x"FF004C34";
      when 4883 => data_o <= x"6F6D75C5";
      when 4884 => data_o <= x"FFFF6576";
      when 4885 => data_o <= x"01FF0006";
      when 4886 => data_o <= x"810012AC";
      when 4887 => data_o <= x"000001DC";
      when 4888 => data_o <= x"FF004C48";
      when 4889 => data_o <= x"6F6D63C5";
      when 4890 => data_o <= x"FFFF6576";
      when 4891 => data_o <= x"01FF000A";
      when 4892 => data_o <= x"890012AC";
      when 4893 => data_o <= x"000001F4";
      when 4894 => data_o <= x"FF004C60";
      when 4895 => data_o <= x"6F6D63C6";
      when 4896 => data_o <= x"FF3E6576";
      when 4897 => data_o <= x"01FF0006";
      when 4898 => data_o <= x"930012AC";
      when 4899 => data_o <= x"0000021C";
      when 4900 => data_o <= x"FF004C78";
      when 4901 => data_o <= x"766F6DC4";
      when 4902 => data_o <= x"FFFFFF65";
      when 4903 => data_o <= x"01FF0006";
      when 4904 => data_o <= x"970012AC";
      when 4905 => data_o <= x"00000234";
      when 4906 => data_o <= x"FF004C90";
      when 4907 => data_o <= x"6C6966C4";
      when 4908 => data_o <= x"FFFFFF6C";
      when 4909 => data_o <= x"01FF000A";
      when 4910 => data_o <= x"A60012AC";
      when 4911 => data_o <= x"0000024C";
      when 4912 => data_o <= x"FF004CA8";
      when 4913 => data_o <= x"617265C5";
      when 4914 => data_o <= x"FFFF6573";
      when 4915 => data_o <= x"01FF0004";
      when 4916 => data_o <= x"B40012AC";
      when 4917 => data_o <= x"00000274";
      when 4918 => data_o <= x"FF004CC0";
      when 4919 => data_o <= x"68736CC6";
      when 4920 => data_o <= x"FF746669";
      when 4921 => data_o <= x"01FF0004";
      when 4922 => data_o <= x"BA0012AC";
      when 4923 => data_o <= x"00000288";
      when 4924 => data_o <= x"FF004CD8";
      when 4925 => data_o <= x"687372C6";
      when 4926 => data_o <= x"FF746669";
      when 4927 => data_o <= x"01FF0003";
      when 4928 => data_o <= x"C10012AC";
      when 4929 => data_o <= x"0000029C";
      when 4930 => data_o <= x"FF004CF0";
      when 4931 => data_o <= x"2A6D75C3";
      when 4932 => data_o <= x"01FF0002";
      when 4933 => data_o <= x"C40012AC";
      when 4934 => data_o <= x"000002A8";
      when 4935 => data_o <= x"FF004D08";
      when 4936 => data_o <= x"FFFF2AC1";
      when 4937 => data_o <= x"01FF0004";
      when 4938 => data_o <= x"C70012AC";
      when 4939 => data_o <= x"000002B0";
      when 4940 => data_o <= x"FF004D1C";
      when 4941 => data_o <= x"2F6D75C6";
      when 4942 => data_o <= x"FF646F6D";
      when 4943 => data_o <= x"01FF000B";
      when 4944 => data_o <= x"ED0012AC";
      when 4945 => data_o <= x"000002C0";
      when 4946 => data_o <= x"FF004D30";
      when 4947 => data_o <= x"2F6D73C6";
      when 4948 => data_o <= x"FF6D6572";
      when 4949 => data_o <= x"01FF000F";
      when 4950 => data_o <= x"F20012AC";
      when 4951 => data_o <= x"000002EC";
      when 4952 => data_o <= x"FF004D48";
      when 4953 => data_o <= x"2F6D66C6";
      when 4954 => data_o <= x"FF646F6D";
      when 4955 => data_o <= x"01FF000B";
      when 4956 => data_o <= x"F90012AC";
      when 4957 => data_o <= x"00000328";
      when 4958 => data_o <= x"FF004D60";
      when 4959 => data_o <= x"6D2F6DC5";
      when 4960 => data_o <= x"FFFF646F";
      when 4961 => data_o <= x"01FF0001";
      when 4962 => data_o <= x"040012AC";
      when 4963 => data_o <= x"01000354";
      when 4964 => data_o <= x"FF004D78";
      when 4965 => data_o <= x"6F6D2FC4";
      when 4966 => data_o <= x"FFFFFF64";
      when 4967 => data_o <= x"01FF0002";
      when 4968 => data_o <= x"050012AC";
      when 4969 => data_o <= x"01000358";
      when 4970 => data_o <= x"FF004D90";
      when 4971 => data_o <= x"646F6DC3";
      when 4972 => data_o <= x"01FF0002";
      when 4973 => data_o <= x"060012AC";
      when 4974 => data_o <= x"01000360";
      when 4975 => data_o <= x"FF004DA8";
      when 4976 => data_o <= x"FFFF2FC1";
      when 4977 => data_o <= x"01FF0003";
      when 4978 => data_o <= x"080012AC";
      when 4979 => data_o <= x"01000368";
      when 4980 => data_o <= x"FF004DBC";
      when 4981 => data_o <= x"6E696DC3";
      when 4982 => data_o <= x"01FF0003";
      when 4983 => data_o <= x"090012AC";
      when 4984 => data_o <= x"01000374";
      when 4985 => data_o <= x"FF004DD0";
      when 4986 => data_o <= x"78616DC3";
      when 4987 => data_o <= x"01FF0003";
      when 4988 => data_o <= x"0A0012AC";
      when 4989 => data_o <= x"01000380";
      when 4990 => data_o <= x"FF004DE4";
      when 4991 => data_o <= x"696D75C4";
      when 4992 => data_o <= x"FFFFFF6E";
      when 4993 => data_o <= x"01FF0003";
      when 4994 => data_o <= x"0B0012AC";
      when 4995 => data_o <= x"0100038C";
      when 4996 => data_o <= x"FF004DF8";
      when 4997 => data_o <= x"616D75C4";
      when 4998 => data_o <= x"FFFFFF78";
      when 4999 => data_o <= x"01FF0002";
      when 5000 => data_o <= x"0D0012AC";
      when 5001 => data_o <= x"01000398";
      when 5002 => data_o <= x"FF004E10";
      when 5003 => data_o <= x"74732FC7";
      when 5004 => data_o <= x"676E6972";
      when 5005 => data_o <= x"01FF0003";
      when 5006 => data_o <= x"0E0012AC";
      when 5007 => data_o <= x"010003A0";
      when 5008 => data_o <= x"FF004E28";
      when 5009 => data_o <= x"746977C6";
      when 5010 => data_o <= x"FF6E6968";
      when 5011 => data_o <= x"01FF0007";
      when 5012 => data_o <= x"0F0012AC";
      when 5013 => data_o <= x"010003AC";
      when 5014 => data_o <= x"FF004E40";
      when 5015 => data_o <= x"FF2A6DC2";
      when 5016 => data_o <= x"01FF0002";
      when 5017 => data_o <= x"140012AC";
      when 5018 => data_o <= x"010003C8";
      when 5019 => data_o <= x"FF004E58";
      when 5020 => data_o <= x"6D2F2AC5";
      when 5021 => data_o <= x"FFFF646F";
      when 5022 => data_o <= x"01FF0002";
      when 5023 => data_o <= x"150012AC";
      when 5024 => data_o <= x"010003D0";
      when 5025 => data_o <= x"FF004E6C";
      when 5026 => data_o <= x"FF2F2AC2";
      when 5027 => data_o <= x"01FF0003";
      when 5028 => data_o <= x"160012AC";
      when 5029 => data_o <= x"010003D8";
      when 5030 => data_o <= x"FF004E84";
      when 5031 => data_o <= x"657962C3";
      when 5032 => data_o <= x"01FF000D";
      when 5033 => data_o <= x"190012AC";
      when 5034 => data_o <= x"010003E4";
      when 5035 => data_o <= x"FF004E98";
      when 5036 => data_o <= x"637263C5";
      when 5037 => data_o <= x"FFFF3233";
      when 5038 => data_o <= x"01FF0008";
      when 5039 => data_o <= x"2A0012AC";
      when 5040 => data_o <= x"01000418";
      when 5041 => data_o <= x"FF004EAC";
      when 5042 => data_o <= x"74616345";
      when 5043 => data_o <= x"FFFF6863";
      when 5044 => data_o <= x"01FF0007";
      when 5045 => data_o <= x"350012AC";
      when 5046 => data_o <= x"01000438";
      when 5047 => data_o <= x"FF004EC4";
      when 5048 => data_o <= x"726874C5";
      when 5049 => data_o <= x"FFFF776F";
      when 5050 => data_o <= x"00FF0001";
      when 5051 => data_o <= x"100012AC";
      when 5052 => data_o <= x"00000454";
      when 5053 => data_o <= x"FF004EDC";
      when 5054 => data_o <= x"756170C5";
      when 5055 => data_o <= x"FFFF6573";
      when 5056 => data_o <= x"00004F48";
      when 5057 => data_o <= x"2F2E2E14";
      when 5058 => data_o <= x"662F2E2E";
      when 5059 => data_o <= x"6874726F";
      when 5060 => data_o <= x"6D69742F";
      when 5061 => data_o <= x"2E676E69";
      when 5062 => data_o <= x"FFFFFF66";
      when 5063 => data_o <= x"02FF0002";
      when 5064 => data_o <= x"010012AC";
      when 5065 => data_o <= x"00000458";
      when 5066 => data_o <= x"FF004EF4";
      when 5067 => data_o <= x"756F63C7";
      when 5068 => data_o <= x"7265746E";
      when 5069 => data_o <= x"02FF0009";
      when 5070 => data_o <= x"040012AC";
      when 5071 => data_o <= x"00000460";
      when 5072 => data_o <= x"FF004F28";
      when 5073 => data_o <= x"FF736DC2";
      when 5074 => data_o <= x"00005304";
      when 5075 => data_o <= x"2F2E2E13";
      when 5076 => data_o <= x"662F2E2E";
      when 5077 => data_o <= x"6874726F";
      when 5078 => data_o <= x"6D756E2F";
      when 5079 => data_o <= x"662E6F69";
      when 5080 => data_o <= x"03FF0003";
      when 5081 => data_o <= x"030012AC";
      when 5082 => data_o <= x"00000484";
      when 5083 => data_o <= x"FF004F40";
      when 5084 => data_o <= x"316F69C4";
      when 5085 => data_o <= x"FFFFFF31";
      when 5086 => data_o <= x"03FF0002";
      when 5087 => data_o <= x"080012AC";
      when 5088 => data_o <= x"00000490";
      when 5089 => data_o <= x"FF004F6C";
      when 5090 => data_o <= x"316F69C4";
      when 5091 => data_o <= x"FFFFFF30";
      when 5092 => data_o <= x"03FF0006";
      when 5093 => data_o <= x"0D0012AC";
      when 5094 => data_o <= x"00000498";
      when 5095 => data_o <= x"FF004F84";
      when 5096 => data_o <= x"726574C9";
      when 5097 => data_o <= x"6D655F6D";
      when 5098 => data_o <= x"FFFF7469";
      when 5099 => data_o <= x"03FF0001";
      when 5100 => data_o <= x"110012AC";
      when 5101 => data_o <= x"000004B0";
      when 5102 => data_o <= x"FF004F9C";
      when 5103 => data_o <= x"707974C4";
      when 5104 => data_o <= x"FFFFFF65";
      when 5105 => data_o <= x"03FF0001";
      when 5106 => data_o <= x"170012AC";
      when 5107 => data_o <= x"000004B4";
      when 5108 => data_o <= x"FF004FB8";
      when 5109 => data_o <= x"797424C5";
      when 5110 => data_o <= x"FFFF6570";
      when 5111 => data_o <= x"000004B8";
      when 5112 => data_o <= x"03FF0000";
      when 5113 => data_o <= x"180012BC";
      when 5114 => data_o <= x"000012B8";
      when 5115 => data_o <= x"FF004FD0";
      when 5116 => data_o <= x"72747309";
      when 5117 => data_o <= x"5F676E69";
      when 5118 => data_o <= x"FFFF7263";
      when 5119 => data_o <= x"000004BB";
      when 5120 => data_o <= x"03FF0000";
      when 5121 => data_o <= x"190012BC";
      when 5122 => data_o <= x"000012B8";
      when 5123 => data_o <= x"FF004FEC";
      when 5124 => data_o <= x"72747309";
      when 5125 => data_o <= x"5F676E69";
      when 5126 => data_o <= x"FFFF6770";
      when 5127 => data_o <= x"03FF0002";
      when 5128 => data_o <= x"1B0012AC";
      when 5129 => data_o <= x"000004C0";
      when 5130 => data_o <= x"FF00500C";
      when 5131 => data_o <= x"726574C7";
      when 5132 => data_o <= x"72635F6D";
      when 5133 => data_o <= x"03FF0002";
      when 5134 => data_o <= x"1C0012AC";
      when 5135 => data_o <= x"000004C8";
      when 5136 => data_o <= x"FF005028";
      when 5137 => data_o <= x"726574C9";
      when 5138 => data_o <= x"61705F6D";
      when 5139 => data_o <= x"FFFF6567";
      when 5140 => data_o <= x"03FF0003";
      when 5141 => data_o <= x"1D0012AC";
      when 5142 => data_o <= x"000004D0";
      when 5143 => data_o <= x"FF005040";
      when 5144 => data_o <= x"726574C9";
      when 5145 => data_o <= x"656B5F6D";
      when 5146 => data_o <= x"FFFF3F79";
      when 5147 => data_o <= x"03FF0005";
      when 5148 => data_o <= x"1E0012AC";
      when 5149 => data_o <= x"000004DC";
      when 5150 => data_o <= x"FF00505C";
      when 5151 => data_o <= x"726574C8";
      when 5152 => data_o <= x"656B5F6D";
      when 5153 => data_o <= x"FFFFFF79";
      when 5154 => data_o <= x"000004F0";
      when 5155 => data_o <= x"03FF0000";
      when 5156 => data_o <= x"2A0012BC";
      when 5157 => data_o <= x"000012B8";
      when 5158 => data_o <= x"FF005078";
      when 5159 => data_o <= x"72657410";
      when 5160 => data_o <= x"65705F6D";
      when 5161 => data_o <= x"6E6F7372";
      when 5162 => data_o <= x"74696C61";
      when 5163 => data_o <= x"FFFFFF79";
      when 5164 => data_o <= x"03FF0003";
      when 5165 => data_o <= x"2C0012AC";
      when 5166 => data_o <= x"00000504";
      when 5167 => data_o <= x"FF005098";
      when 5168 => data_o <= x"3D6F69C7";
      when 5169 => data_o <= x"6D726574";
      when 5170 => data_o <= x"03FF0002";
      when 5171 => data_o <= x"2F0012AC";
      when 5172 => data_o <= x"00000510";
      when 5173 => data_o <= x"FF0050BC";
      when 5174 => data_o <= x"726570D0";
      when 5175 => data_o <= x"616E6F73";
      when 5176 => data_o <= x"7974696C";
      when 5177 => data_o <= x"6578655F";
      when 5178 => data_o <= x"FFFFFF63";
      when 5179 => data_o <= x"03FF0002";
      when 5180 => data_o <= x"330012AC";
      when 5181 => data_o <= x"00000518";
      when 5182 => data_o <= x"FF0050D4";
      when 5183 => data_o <= x"696D65C4";
      when 5184 => data_o <= x"FFFFFF74";
      when 5185 => data_o <= x"03FF0002";
      when 5186 => data_o <= x"340012AC";
      when 5187 => data_o <= x"00000520";
      when 5188 => data_o <= x"FF0050F8";
      when 5189 => data_o <= x"FF7263C2";
      when 5190 => data_o <= x"03FF0002";
      when 5191 => data_o <= x"350012AC";
      when 5192 => data_o <= x"00000528";
      when 5193 => data_o <= x"FF005110";
      when 5194 => data_o <= x"676170C4";
      when 5195 => data_o <= x"FFFFFF65";
      when 5196 => data_o <= x"03FF0002";
      when 5197 => data_o <= x"360012AC";
      when 5198 => data_o <= x"00000530";
      when 5199 => data_o <= x"FF005124";
      when 5200 => data_o <= x"79656BC4";
      when 5201 => data_o <= x"FFFFFF3F";
      when 5202 => data_o <= x"03FF0002";
      when 5203 => data_o <= x"370012AC";
      when 5204 => data_o <= x"00000538";
      when 5205 => data_o <= x"FF00513C";
      when 5206 => data_o <= x"79656BC3";
      when 5207 => data_o <= x"03FF0002";
      when 5208 => data_o <= x"3F0012AC";
      when 5209 => data_o <= x"00000558";
      when 5210 => data_o <= x"FF005154";
      when 5211 => data_o <= x"617073C5";
      when 5212 => data_o <= x"FFFF6563";
      when 5213 => data_o <= x"03FF0005";
      when 5214 => data_o <= x"400012AC";
      when 5215 => data_o <= x"00000560";
      when 5216 => data_o <= x"FF005168";
      when 5217 => data_o <= x"617073C6";
      when 5218 => data_o <= x"FF736563";
      when 5219 => data_o <= x"03FF0004";
      when 5220 => data_o <= x"470012AC";
      when 5221 => data_o <= x"00000574";
      when 5222 => data_o <= x"FF005180";
      when 5223 => data_o <= x"676964C5";
      when 5224 => data_o <= x"FFFF7469";
      when 5225 => data_o <= x"03FF0003";
      when 5226 => data_o <= x"480012AC";
      when 5227 => data_o <= x"00000584";
      when 5228 => data_o <= x"FF005198";
      when 5229 => data_o <= x"FF233CC2";
      when 5230 => data_o <= x"03FF0004";
      when 5231 => data_o <= x"4A0012AC";
      when 5232 => data_o <= x"00000590";
      when 5233 => data_o <= x"FF0051B0";
      when 5234 => data_o <= x"6C6F68C4";
      when 5235 => data_o <= x"FFFFFF64";
      when 5236 => data_o <= x"03FF000D";
      when 5237 => data_o <= x"4C0012AC";
      when 5238 => data_o <= x"000005A0";
      when 5239 => data_o <= x"FF0051C4";
      when 5240 => data_o <= x"FFFF23C1";
      when 5241 => data_o <= x"03FF0004";
      when 5242 => data_o <= x"540012AC";
      when 5243 => data_o <= x"000005D4";
      when 5244 => data_o <= x"FF0051DC";
      when 5245 => data_o <= x"FF7323C2";
      when 5246 => data_o <= x"03FF0004";
      when 5247 => data_o <= x"550012AC";
      when 5248 => data_o <= x"000005E4";
      when 5249 => data_o <= x"FF0051F0";
      when 5250 => data_o <= x"676973C4";
      when 5251 => data_o <= x"FFFFFF6E";
      when 5252 => data_o <= x"03FF0003";
      when 5253 => data_o <= x"560012AC";
      when 5254 => data_o <= x"000005F4";
      when 5255 => data_o <= x"FF005204";
      when 5256 => data_o <= x"FF3E23C2";
      when 5257 => data_o <= x"03FF0003";
      when 5258 => data_o <= x"570012AC";
      when 5259 => data_o <= x"00000600";
      when 5260 => data_o <= x"FF00521C";
      when 5261 => data_o <= x"722E73C3";
      when 5262 => data_o <= x"03FF0006";
      when 5263 => data_o <= x"580012AC";
      when 5264 => data_o <= x"0000060C";
      when 5265 => data_o <= x"FF005230";
      when 5266 => data_o <= x"722E64C3";
      when 5267 => data_o <= x"03FF0002";
      when 5268 => data_o <= x"5A0012AC";
      when 5269 => data_o <= x"00000624";
      when 5270 => data_o <= x"FF005244";
      when 5271 => data_o <= x"722E75C3";
      when 5272 => data_o <= x"03FF0002";
      when 5273 => data_o <= x"5B0012AC";
      when 5274 => data_o <= x"0000062C";
      when 5275 => data_o <= x"FF005258";
      when 5276 => data_o <= x"FF722EC2";
      when 5277 => data_o <= x"03FF0003";
      when 5278 => data_o <= x"5C0012AC";
      when 5279 => data_o <= x"00000634";
      when 5280 => data_o <= x"FF00526C";
      when 5281 => data_o <= x"FF2E64C2";
      when 5282 => data_o <= x"03FF0002";
      when 5283 => data_o <= x"5D0012AC";
      when 5284 => data_o <= x"00000640";
      when 5285 => data_o <= x"FF005280";
      when 5286 => data_o <= x"FF2E75C2";
      when 5287 => data_o <= x"03FF0006";
      when 5288 => data_o <= x"5E0012AC";
      when 5289 => data_o <= x"00000648";
      when 5290 => data_o <= x"FF005294";
      when 5291 => data_o <= x"FFFF2EC1";
      when 5292 => data_o <= x"03FF0001";
      when 5293 => data_o <= x"610012AC";
      when 5294 => data_o <= x"00000660";
      when 5295 => data_o <= x"FF0052A8";
      when 5296 => data_o <= x"FFFF3FC1";
      when 5297 => data_o <= x"03FF0007";
      when 5298 => data_o <= x"620012AC";
      when 5299 => data_o <= x"00000664";
      when 5300 => data_o <= x"FF0052BC";
      when 5301 => data_o <= x"3E233CC3";
      when 5302 => data_o <= x"03FF0008";
      when 5303 => data_o <= x"630012AC";
      when 5304 => data_o <= x"00000680";
      when 5305 => data_o <= x"FF0052D0";
      when 5306 => data_o <= x"782E68C3";
      when 5307 => data_o <= x"03FF0026";
      when 5308 => data_o <= x"680012AC";
      when 5309 => data_o <= x"000006A0";
      when 5310 => data_o <= x"FF0052E4";
      when 5311 => data_o <= x"636361C6";
      when 5312 => data_o <= x"FF747065";
      when 5313 => data_o <= x"00005448";
      when 5314 => data_o <= x"2F2E2E13";
      when 5315 => data_o <= x"662F2E2E";
      when 5316 => data_o <= x"6874726F";
      when 5317 => data_o <= x"616C662F";
      when 5318 => data_o <= x"662E6873";
      when 5319 => data_o <= x"04FF0005";
      when 5320 => data_o <= x"090012AC";
      when 5321 => data_o <= x"0000073C";
      when 5322 => data_o <= x"FF0052F8";
      when 5323 => data_o <= x"495053C7";
      when 5324 => data_o <= x"72656678";
      when 5325 => data_o <= x"04FF000B";
      when 5326 => data_o <= x"0E0012AC";
      when 5327 => data_o <= x"00000750";
      when 5328 => data_o <= x"FF005328";
      when 5329 => data_o <= x"495053CA";
      when 5330 => data_o <= x"72646461";
      when 5331 => data_o <= x"FF737365";
      when 5332 => data_o <= x"04FF0004";
      when 5333 => data_o <= x"190012AC";
      when 5334 => data_o <= x"0000077C";
      when 5335 => data_o <= x"FF005340";
      when 5336 => data_o <= x"495053C5";
      when 5337 => data_o <= x"FFFF5253";
      when 5338 => data_o <= x"04FF0005";
      when 5339 => data_o <= x"1D0012AC";
      when 5340 => data_o <= x"0000078C";
      when 5341 => data_o <= x"FF00535C";
      when 5342 => data_o <= x"495053C7";
      when 5343 => data_o <= x"74696177";
      when 5344 => data_o <= x"04FF0005";
      when 5345 => data_o <= x"200012AC";
      when 5346 => data_o <= x"000007A0";
      when 5347 => data_o <= x"FF005374";
      when 5348 => data_o <= x"495053C5";
      when 5349 => data_o <= x"FFFF4449";
      when 5350 => data_o <= x"04FF0008";
      when 5351 => data_o <= x"260012AC";
      when 5352 => data_o <= x"000007B4";
      when 5353 => data_o <= x"FF00538C";
      when 5354 => data_o <= x"495053CA";
      when 5355 => data_o <= x"73617265";
      when 5356 => data_o <= x"FF4B3465";
      when 5357 => data_o <= x"04FF0003";
      when 5358 => data_o <= x"2C0012AC";
      when 5359 => data_o <= x"000007D4";
      when 5360 => data_o <= x"FF0053A4";
      when 5361 => data_o <= x"495053C7";
      when 5362 => data_o <= x"65747962";
      when 5363 => data_o <= x"04FF0011";
      when 5364 => data_o <= x"310012AC";
      when 5365 => data_o <= x"000007E0";
      when 5366 => data_o <= x"FF0053C0";
      when 5367 => data_o <= x"50535FC8";
      when 5368 => data_o <= x"766F6D49";
      when 5369 => data_o <= x"FFFFFF65";
      when 5370 => data_o <= x"04FF0016";
      when 5371 => data_o <= x"430012AC";
      when 5372 => data_o <= x"00000824";
      when 5373 => data_o <= x"FF0053D8";
      when 5374 => data_o <= x"495053C7";
      when 5375 => data_o <= x"74736574";
      when 5376 => data_o <= x"04FF000B";
      when 5377 => data_o <= x"530012AC";
      when 5378 => data_o <= x"0000087C";
      when 5379 => data_o <= x"FF0053F4";
      when 5380 => data_o <= x"495053C7";
      when 5381 => data_o <= x"65766F6D";
      when 5382 => data_o <= x"04FF0005";
      when 5383 => data_o <= x"5D0012AC";
      when 5384 => data_o <= x"000008A8";
      when 5385 => data_o <= x"FF00540C";
      when 5386 => data_o <= x"495053C4";
      when 5387 => data_o <= x"FFFFFF21";
      when 5388 => data_o <= x"04FF000D";
      when 5389 => data_o <= x"630012AC";
      when 5390 => data_o <= x"000008BC";
      when 5391 => data_o <= x"FF005424";
      when 5392 => data_o <= x"495053C4";
      when 5393 => data_o <= x"FFFFFF40";
      when 5394 => data_o <= x"000055F4";
      when 5395 => data_o <= x"2F2E2E13";
      when 5396 => data_o <= x"662F2E2E";
      when 5397 => data_o <= x"6874726F";
      when 5398 => data_o <= x"6D6F632F";
      when 5399 => data_o <= x"662E616D";
      when 5400 => data_o <= x"05FF0004";
      when 5401 => data_o <= x"220012AC";
      when 5402 => data_o <= x"000008F0";
      when 5403 => data_o <= x"FF00543C";
      when 5404 => data_o <= x"4D4F52C4";
      when 5405 => data_o <= x"FFFFFF21";
      when 5406 => data_o <= x"05FF000D";
      when 5407 => data_o <= x"260012AC";
      when 5408 => data_o <= x"00000900";
      when 5409 => data_o <= x"FF00546C";
      when 5410 => data_o <= x"4D4F52C5";
      when 5411 => data_o <= x"FFFF2143";
      when 5412 => data_o <= x"05FF000A";
      when 5413 => data_o <= x"2F0012AC";
      when 5414 => data_o <= x"00000934";
      when 5415 => data_o <= x"FF005484";
      when 5416 => data_o <= x"4D4F52C7";
      when 5417 => data_o <= x"65766F6D";
      when 5418 => data_o <= x"05FF0003";
      when 5419 => data_o <= x"3E0012AC";
      when 5420 => data_o <= x"0000095C";
      when 5421 => data_o <= x"FF00549C";
      when 5422 => data_o <= x"6D6172C3";
      when 5423 => data_o <= x"05FF0003";
      when 5424 => data_o <= x"3F0012AC";
      when 5425 => data_o <= x"00000968";
      when 5426 => data_o <= x"FF0054B4";
      when 5427 => data_o <= x"6D6F72C3";
      when 5428 => data_o <= x"05FF0007";
      when 5429 => data_o <= x"400012AC";
      when 5430 => data_o <= x"00000974";
      when 5431 => data_o <= x"FF0054C8";
      when 5432 => data_o <= x"FFFF68C1";
      when 5433 => data_o <= x"05FF0004";
      when 5434 => data_o <= x"410012AC";
      when 5435 => data_o <= x"00000990";
      when 5436 => data_o <= x"FF0054DC";
      when 5437 => data_o <= x"FF782CC2";
      when 5438 => data_o <= x"05FF0002";
      when 5439 => data_o <= x"420012AC";
      when 5440 => data_o <= x"000009A0";
      when 5441 => data_o <= x"FF0054F0";
      when 5442 => data_o <= x"FF632CC2";
      when 5443 => data_o <= x"05FF0002";
      when 5444 => data_o <= x"430012AC";
      when 5445 => data_o <= x"000009A8";
      when 5446 => data_o <= x"FF005504";
      when 5447 => data_o <= x"FF682CC2";
      when 5448 => data_o <= x"05FF0004";
      when 5449 => data_o <= x"440012AC";
      when 5450 => data_o <= x"000009B0";
      when 5451 => data_o <= x"FF005518";
      when 5452 => data_o <= x"FF642CC2";
      when 5453 => data_o <= x"05FF0005";
      when 5454 => data_o <= x"450012AC";
      when 5455 => data_o <= x"000009C0";
      when 5456 => data_o <= x"FF00552C";
      when 5457 => data_o <= x"FFFF2CC1";
      when 5458 => data_o <= x"05FF0004";
      when 5459 => data_o <= x"470012AC";
      when 5460 => data_o <= x"000009D4";
      when 5461 => data_o <= x"FF005540";
      when 5462 => data_o <= x"782C63C3";
      when 5463 => data_o <= x"05FF0002";
      when 5464 => data_o <= x"4A0012AC";
      when 5465 => data_o <= x"000009E4";
      when 5466 => data_o <= x"FF005554";
      when 5467 => data_o <= x"632C63C3";
      when 5468 => data_o <= x"05FF0002";
      when 5469 => data_o <= x"4B0012AC";
      when 5470 => data_o <= x"000009EC";
      when 5471 => data_o <= x"FF005568";
      when 5472 => data_o <= x"682C63C3";
      when 5473 => data_o <= x"05FF0004";
      when 5474 => data_o <= x"4C0012AC";
      when 5475 => data_o <= x"000009F4";
      when 5476 => data_o <= x"FF00557C";
      when 5477 => data_o <= x"642C63C3";
      when 5478 => data_o <= x"05FF0005";
      when 5479 => data_o <= x"4D0012AC";
      when 5480 => data_o <= x"00000A04";
      when 5481 => data_o <= x"FF005590";
      when 5482 => data_o <= x"FF2C63C2";
      when 5483 => data_o <= x"05FF0002";
      when 5484 => data_o <= x"520012AC";
      when 5485 => data_o <= x"00000A18";
      when 5486 => data_o <= x"FF0055A4";
      when 5487 => data_o <= x"6E6F63C4";
      when 5488 => data_o <= x"FFFFFF74";
      when 5489 => data_o <= x"05FF000E";
      when 5490 => data_o <= x"550012AC";
      when 5491 => data_o <= x"00000A20";
      when 5492 => data_o <= x"FF0055B8";
      when 5493 => data_o <= x"64695FC7";
      when 5494 => data_o <= x"2C617461";
      when 5495 => data_o <= x"05FF000F";
      when 5496 => data_o <= x"5B0012AC";
      when 5497 => data_o <= x"00000A58";
      when 5498 => data_o <= x"FF0055D0";
      when 5499 => data_o <= x"616469C6";
      when 5500 => data_o <= x"FF2C6174";
      when 5501 => data_o <= x"000059B8";
      when 5502 => data_o <= x"2F2E2E15";
      when 5503 => data_o <= x"662F2E2E";
      when 5504 => data_o <= x"6874726F";
      when 5505 => data_o <= x"6D6F632F";
      when 5506 => data_o <= x"656C6970";
      when 5507 => data_o <= x"FFFF662E";
      when 5508 => data_o <= x"FFFFF214";
      when 5509 => data_o <= x"06FF0000";
      when 5510 => data_o <= x"060012BC";
      when 5511 => data_o <= x"000012B8";
      when 5512 => data_o <= x"FF0055E8";
      when 5513 => data_o <= x"6E616807";
      when 5514 => data_o <= x"72656C64";
      when 5515 => data_o <= x"FFFFF218";
      when 5516 => data_o <= x"06FF0000";
      when 5517 => data_o <= x"070012BC";
      when 5518 => data_o <= x"000012B8";
      when 5519 => data_o <= x"FF005620";
      when 5520 => data_o <= x"73616204";
      when 5521 => data_o <= x"FFFFFF65";
      when 5522 => data_o <= x"FFFFF21C";
      when 5523 => data_o <= x"06FF0000";
      when 5524 => data_o <= x"080012BC";
      when 5525 => data_o <= x"000012B8";
      when 5526 => data_o <= x"FF00563C";
      when 5527 => data_o <= x"FF706802";
      when 5528 => data_o <= x"FFFFF220";
      when 5529 => data_o <= x"06FF0000";
      when 5530 => data_o <= x"090012BC";
      when 5531 => data_o <= x"000012B8";
      when 5532 => data_o <= x"FF005658";
      when 5533 => data_o <= x"FF706302";
      when 5534 => data_o <= x"FFFFF224";
      when 5535 => data_o <= x"06FF0000";
      when 5536 => data_o <= x"0A0012BC";
      when 5537 => data_o <= x"000012B8";
      when 5538 => data_o <= x"FF005670";
      when 5539 => data_o <= x"FF706402";
      when 5540 => data_o <= x"FFFFF228";
      when 5541 => data_o <= x"06FF0000";
      when 5542 => data_o <= x"0B0012BC";
      when 5543 => data_o <= x"000012B8";
      when 5544 => data_o <= x"FF005688";
      when 5545 => data_o <= x"61747305";
      when 5546 => data_o <= x"FFFF6574";
      when 5547 => data_o <= x"FFFFF22C";
      when 5548 => data_o <= x"06FF0000";
      when 5549 => data_o <= x"0C0012BC";
      when 5550 => data_o <= x"000012B8";
      when 5551 => data_o <= x"FF0056A0";
      when 5552 => data_o <= x"72756307";
      when 5553 => data_o <= x"746E6572";
      when 5554 => data_o <= x"FFFFF234";
      when 5555 => data_o <= x"06FF0000";
      when 5556 => data_o <= x"0D0012BC";
      when 5557 => data_o <= x"000012B8";
      when 5558 => data_o <= x"FF0056BC";
      when 5559 => data_o <= x"756F7309";
      when 5560 => data_o <= x"2D656372";
      when 5561 => data_o <= x"FFFF6469";
      when 5562 => data_o <= x"FFFFF230";
      when 5563 => data_o <= x"06FF0000";
      when 5564 => data_o <= x"0E0012BC";
      when 5565 => data_o <= x"000012B8";
      when 5566 => data_o <= x"FF0056D8";
      when 5567 => data_o <= x"7265700B";
      when 5568 => data_o <= x"616E6F73";
      when 5569 => data_o <= x"7974696C";
      when 5570 => data_o <= x"FFFFF238";
      when 5571 => data_o <= x"06FF0000";
      when 5572 => data_o <= x"0F0012BC";
      when 5573 => data_o <= x"000012B8";
      when 5574 => data_o <= x"FF0056F8";
      when 5575 => data_o <= x"62697404";
      when 5576 => data_o <= x"FFFFFF73";
      when 5577 => data_o <= x"FFFFF23C";
      when 5578 => data_o <= x"06FF0000";
      when 5579 => data_o <= x"100012BC";
      when 5580 => data_o <= x"000012B8";
      when 5581 => data_o <= x"FF005718";
      when 5582 => data_o <= x"62697404";
      when 5583 => data_o <= x"FFFFFF62";
      when 5584 => data_o <= x"FFFFF240";
      when 5585 => data_o <= x"06FF0000";
      when 5586 => data_o <= x"110012BC";
      when 5587 => data_o <= x"000012B8";
      when 5588 => data_o <= x"FF005734";
      when 5589 => data_o <= x"6E693E03";
      when 5590 => data_o <= x"FFFFF248";
      when 5591 => data_o <= x"06FF0000";
      when 5592 => data_o <= x"120012BC";
      when 5593 => data_o <= x"000012B8";
      when 5594 => data_o <= x"FF005750";
      when 5595 => data_o <= x"775F6306";
      when 5596 => data_o <= x"FF736469";
      when 5597 => data_o <= x"FFFFF24D";
      when 5598 => data_o <= x"06FF0000";
      when 5599 => data_o <= x"130012BC";
      when 5600 => data_o <= x"000012B8";
      when 5601 => data_o <= x"FF005768";
      when 5602 => data_o <= x"635F630A";
      when 5603 => data_o <= x"73657361";
      when 5604 => data_o <= x"FF736E65";
      when 5605 => data_o <= x"FFFFF264";
      when 5606 => data_o <= x"06FF0000";
      when 5607 => data_o <= x"150012BC";
      when 5608 => data_o <= x"000012B8";
      when 5609 => data_o <= x"FF005784";
      when 5610 => data_o <= x"6E6F6307";
      when 5611 => data_o <= x"74786574";
      when 5612 => data_o <= x"FFFFF334";
      when 5613 => data_o <= x"06FF0000";
      when 5614 => data_o <= x"160012BC";
      when 5615 => data_o <= x"000012B8";
      when 5616 => data_o <= x"FF0057A4";
      when 5617 => data_o <= x"726F660E";
      when 5618 => data_o <= x"772D6874";
      when 5619 => data_o <= x"6C64726F";
      when 5620 => data_o <= x"FF747369";
      when 5621 => data_o <= x"FFFFF268";
      when 5622 => data_o <= x"06FF0000";
      when 5623 => data_o <= x"170012BC";
      when 5624 => data_o <= x"000012B8";
      when 5625 => data_o <= x"FF0057C0";
      when 5626 => data_o <= x"646C6803";
      when 5627 => data_o <= x"FFFFF244";
      when 5628 => data_o <= x"06FF0000";
      when 5629 => data_o <= x"180012BC";
      when 5630 => data_o <= x"000012B8";
      when 5631 => data_o <= x"FF0057E4";
      when 5632 => data_o <= x"6B6C6203";
      when 5633 => data_o <= x"FFFFF26C";
      when 5634 => data_o <= x"06FF0000";
      when 5635 => data_o <= x"190012BC";
      when 5636 => data_o <= x"000012B8";
      when 5637 => data_o <= x"FF0057FC";
      when 5638 => data_o <= x"62697403";
      when 5639 => data_o <= x"00000040";
      when 5640 => data_o <= x"06FF0000";
      when 5641 => data_o <= x"1B0012BC";
      when 5642 => data_o <= x"000012B8";
      when 5643 => data_o <= x"FF005814";
      when 5644 => data_o <= x"61707C05";
      when 5645 => data_o <= x"FFFF7C64";
      when 5646 => data_o <= x"FFFFF2F4";
      when 5647 => data_o <= x"06FF0000";
      when 5648 => data_o <= x"1C0012BC";
      when 5649 => data_o <= x"000012B8";
      when 5650 => data_o <= x"FF00582C";
      when 5651 => data_o <= x"64617003";
      when 5652 => data_o <= x"00001000";
      when 5653 => data_o <= x"06FF0000";
      when 5654 => data_o <= x"1D0012BC";
      when 5655 => data_o <= x"000012B8";
      when 5656 => data_o <= x"FF005848";
      when 5657 => data_o <= x"4D415207";
      when 5658 => data_o <= x"657A6973";
      when 5659 => data_o <= x"00008000";
      when 5660 => data_o <= x"06FF0000";
      when 5661 => data_o <= x"1E0012BC";
      when 5662 => data_o <= x"000012B8";
      when 5663 => data_o <= x"FF005860";
      when 5664 => data_o <= x"4D4F5207";
      when 5665 => data_o <= x"657A6973";
      when 5666 => data_o <= x"00000100";
      when 5667 => data_o <= x"06FF0000";
      when 5668 => data_o <= x"1F0012BC";
      when 5669 => data_o <= x"000012B8";
      when 5670 => data_o <= x"FF00587C";
      when 5671 => data_o <= x"4950530E";
      when 5672 => data_o <= x"73616C66";
      when 5673 => data_o <= x"6F6C4268";
      when 5674 => data_o <= x"FF736B63";
      when 5675 => data_o <= x"06FF0001";
      when 5676 => data_o <= x"240012AC";
      when 5677 => data_o <= x"00000A94";
      when 5678 => data_o <= x"FF005898";
      when 5679 => data_o <= x"756C46C8";
      when 5680 => data_o <= x"694C6873";
      when 5681 => data_o <= x"FFFFFF74";
      when 5682 => data_o <= x"06FF0001";
      when 5683 => data_o <= x"250012AC";
      when 5684 => data_o <= x"00000A98";
      when 5685 => data_o <= x"FF0058B8";
      when 5686 => data_o <= x"77654EC8";
      when 5687 => data_o <= x"756F7247";
      when 5688 => data_o <= x"FFFFFF70";
      when 5689 => data_o <= x"06FF0007";
      when 5690 => data_o <= x"270012AC";
      when 5691 => data_o <= x"00000A9C";
      when 5692 => data_o <= x"FF0058D4";
      when 5693 => data_o <= x"656C43C7";
      when 5694 => data_o <= x"52497261";
      when 5695 => data_o <= x"06FF0006";
      when 5696 => data_o <= x"2A0012AC";
      when 5697 => data_o <= x"00000AB8";
      when 5698 => data_o <= x"FF0058F0";
      when 5699 => data_o <= x"707041C8";
      when 5700 => data_o <= x"49646E65";
      when 5701 => data_o <= x"FFFFFF52";
      when 5702 => data_o <= x"06FF0011";
      when 5703 => data_o <= x"2F0012AC";
      when 5704 => data_o <= x"00000AD0";
      when 5705 => data_o <= x"FF005908";
      when 5706 => data_o <= x"706D49C8";
      when 5707 => data_o <= x"6963696C";
      when 5708 => data_o <= x"FFFFFF74";
      when 5709 => data_o <= x"06FF0014";
      when 5710 => data_o <= x"3C0012AC";
      when 5711 => data_o <= x"00000B14";
      when 5712 => data_o <= x"FF005924";
      when 5713 => data_o <= x"707845C8";
      when 5714 => data_o <= x"6963696C";
      when 5715 => data_o <= x"FFFFFF74";
      when 5716 => data_o <= x"06FF0013";
      when 5717 => data_o <= x"480012AC";
      when 5718 => data_o <= x"00000B64";
      when 5719 => data_o <= x"FF005940";
      when 5720 => data_o <= x"726148C7";
      when 5721 => data_o <= x"74694C64";
      when 5722 => data_o <= x"06FF0009";
      when 5723 => data_o <= x"690012AC";
      when 5724 => data_o <= x"00000C08";
      when 5725 => data_o <= x"FF00595C";
      when 5726 => data_o <= x"74696CC8";
      when 5727 => data_o <= x"6C617265";
      when 5728 => data_o <= x"FFFFFF2C";
      when 5729 => data_o <= x"06FF0007";
      when 5730 => data_o <= x"6F0012AC";
      when 5731 => data_o <= x"00000C2C";
      when 5732 => data_o <= x"FF005974";
      when 5733 => data_o <= x"6D6F63C8";
      when 5734 => data_o <= x"656C6970";
      when 5735 => data_o <= x"FFFFFF2C";
      when 5736 => data_o <= x"06FF0010";
      when 5737 => data_o <= x"730012AC";
      when 5738 => data_o <= x"00000C48";
      when 5739 => data_o <= x"FF005990";
      when 5740 => data_o <= x"78652CC5";
      when 5741 => data_o <= x"FFFF7469";
      when 5742 => data_o <= x"00005C18";
      when 5743 => data_o <= x"2F2E2E13";
      when 5744 => data_o <= x"662F2E2E";
      when 5745 => data_o <= x"6874726F";
      when 5746 => data_o <= x"6F6F742F";
      when 5747 => data_o <= x"662E736C";
      when 5748 => data_o <= x"07FF0008";
      when 5749 => data_o <= x"030012AC";
      when 5750 => data_o <= x"00000C88";
      when 5751 => data_o <= x"FF0059AC";
      when 5752 => data_o <= x"FF2E3BC2";
      when 5753 => data_o <= x"07FF0003";
      when 5754 => data_o <= x"070012AC";
      when 5755 => data_o <= x"00000CA8";
      when 5756 => data_o <= x"FF0059DC";
      when 5757 => data_o <= x"6C6F6348";
      when 5758 => data_o <= x"7A69726F";
      when 5759 => data_o <= x"FFFFFF65";
      when 5760 => data_o <= x"07FF0003";
      when 5761 => data_o <= x"0A0012AC";
      when 5762 => data_o <= x"00000CB4";
      when 5763 => data_o <= x"FF0059F0";
      when 5764 => data_o <= x"656874CA";
      when 5765 => data_o <= x"6D3D656D";
      when 5766 => data_o <= x"FF6F6E6F";
      when 5767 => data_o <= x"07FF0003";
      when 5768 => data_o <= x"0B0012AC";
      when 5769 => data_o <= x"00000CC0";
      when 5770 => data_o <= x"FF005A0C";
      when 5771 => data_o <= x"656874CB";
      when 5772 => data_o <= x"633D656D";
      when 5773 => data_o <= x"726F6C6F";
      when 5774 => data_o <= x"07FF0005";
      when 5775 => data_o <= x"0E0012AC";
      when 5776 => data_o <= x"00000CCC";
      when 5777 => data_o <= x"FF005A28";
      when 5778 => data_o <= x"637365C4";
      when 5779 => data_o <= x"FFFFFF5B";
      when 5780 => data_o <= x"07FF0002";
      when 5781 => data_o <= x"0F0012AC";
      when 5782 => data_o <= x"00000CE0";
      when 5783 => data_o <= x"FF005A44";
      when 5784 => data_o <= x"637365C5";
      when 5785 => data_o <= x"FFFF305B";
      when 5786 => data_o <= x"07FF0002";
      when 5787 => data_o <= x"100012AC";
      when 5788 => data_o <= x"00000CE8";
      when 5789 => data_o <= x"FF005A5C";
      when 5790 => data_o <= x"637365C5";
      when 5791 => data_o <= x"FFFF315B";
      when 5792 => data_o <= x"07FF0002";
      when 5793 => data_o <= x"110012AC";
      when 5794 => data_o <= x"00000CF0";
      when 5795 => data_o <= x"FF005A74";
      when 5796 => data_o <= x"FF6D5DC2";
      when 5797 => data_o <= x"07FF0003";
      when 5798 => data_o <= x"130012AC";
      when 5799 => data_o <= x"00000CF8";
      when 5800 => data_o <= x"FF005A8C";
      when 5801 => data_o <= x"6C6F43C9";
      when 5802 => data_o <= x"6F4E726F";
      when 5803 => data_o <= x"FFFF656E";
      when 5804 => data_o <= x"07FF0003";
      when 5805 => data_o <= x"140012AC";
      when 5806 => data_o <= x"00000D04";
      when 5807 => data_o <= x"FF005AA0";
      when 5808 => data_o <= x"6C6F63C7";
      when 5809 => data_o <= x"785F726F";
      when 5810 => data_o <= x"07FF0003";
      when 5811 => data_o <= x"150012AC";
      when 5812 => data_o <= x"00000D10";
      when 5813 => data_o <= x"FF005ABC";
      when 5814 => data_o <= x"6C6F63C8";
      when 5815 => data_o <= x"785F726F";
      when 5816 => data_o <= x"FFFFFF64";
      when 5817 => data_o <= x"07FF0003";
      when 5818 => data_o <= x"160012AC";
      when 5819 => data_o <= x"00000D1C";
      when 5820 => data_o <= x"FF005AD4";
      when 5821 => data_o <= x"6C6F43C7";
      when 5822 => data_o <= x"6948726F";
      when 5823 => data_o <= x"07FF0003";
      when 5824 => data_o <= x"170012AC";
      when 5825 => data_o <= x"00000D28";
      when 5826 => data_o <= x"FF005AF0";
      when 5827 => data_o <= x"6C6F43C8";
      when 5828 => data_o <= x"6544726F";
      when 5829 => data_o <= x"FFFFFF66";
      when 5830 => data_o <= x"07FF0003";
      when 5831 => data_o <= x"180012AC";
      when 5832 => data_o <= x"00000D34";
      when 5833 => data_o <= x"FF005B08";
      when 5834 => data_o <= x"6C6F43C9";
      when 5835 => data_o <= x"6F43726F";
      when 5836 => data_o <= x"FFFF706D";
      when 5837 => data_o <= x"07FF0003";
      when 5838 => data_o <= x"190012AC";
      when 5839 => data_o <= x"00000D40";
      when 5840 => data_o <= x"FF005B24";
      when 5841 => data_o <= x"6C6F43C8";
      when 5842 => data_o <= x"6D49726F";
      when 5843 => data_o <= x"FFFFFF6D";
      when 5844 => data_o <= x"07FF0003";
      when 5845 => data_o <= x"1A0012AC";
      when 5846 => data_o <= x"00000D4C";
      when 5847 => data_o <= x"FF005B40";
      when 5848 => data_o <= x"6C6F43C9";
      when 5849 => data_o <= x"6D49726F";
      when 5850 => data_o <= x"FFFF416D";
      when 5851 => data_o <= x"07FF0001";
      when 5852 => data_o <= x"1B0012AC";
      when 5853 => data_o <= x"00000D58";
      when 5854 => data_o <= x"FF005B5C";
      when 5855 => data_o <= x"6C6F43CA";
      when 5856 => data_o <= x"704F726F";
      when 5857 => data_o <= x"FF646F63";
      when 5858 => data_o <= x"00000D5C";
      when 5859 => data_o <= x"07FF0000";
      when 5860 => data_o <= x"300012BC";
      when 5861 => data_o <= x"000012B8";
      when 5862 => data_o <= x"FF005B78";
      when 5863 => data_o <= x"726F770A";
      when 5864 => data_o <= x"6C6F6364";
      when 5865 => data_o <= x"FF73726F";
      when 5866 => data_o <= x"07FF000D";
      when 5867 => data_o <= x"330012AC";
      when 5868 => data_o <= x"00000D6C";
      when 5869 => data_o <= x"FF005B98";
      when 5870 => data_o <= x"6C6F43C9";
      when 5871 => data_o <= x"6F57726F";
      when 5872 => data_o <= x"FFFF6472";
      when 5873 => data_o <= x"07FF000D";
      when 5874 => data_o <= x"490012AC";
      when 5875 => data_o <= x"00000DA0";
      when 5876 => data_o <= x"FF005BB4";
      when 5877 => data_o <= x"FF732EC2";
      when 5878 => data_o <= x"07FF0026";
      when 5879 => data_o <= x"530012AC";
      when 5880 => data_o <= x"00000DD4";
      when 5881 => data_o <= x"FF005BD0";
      when 5882 => data_o <= x"6D7564C4";
      when 5883 => data_o <= x"FFFFFF70";
      when 5884 => data_o <= x"07FF0006";
      when 5885 => data_o <= x"6A0012AC";
      when 5886 => data_o <= x"00000E6C";
      when 5887 => data_o <= x"FF005BE4";
      when 5888 => data_o <= x"523E4E43";
      when 5889 => data_o <= x"07FF0006";
      when 5890 => data_o <= x"770012AC";
      when 5891 => data_o <= x"00000E84";
      when 5892 => data_o <= x"FF005BFC";
      when 5893 => data_o <= x"3E524E43";
      when 5894 => data_o <= x"00005EC0";
      when 5895 => data_o <= x"2F2E2E17";
      when 5896 => data_o <= x"662F2E2E";
      when 5897 => data_o <= x"6874726F";
      when 5898 => data_o <= x"746E692F";
      when 5899 => data_o <= x"72707265";
      when 5900 => data_o <= x"662E7465";
      when 5901 => data_o <= x"08FF0005";
      when 5902 => data_o <= x"040012AC";
      when 5903 => data_o <= x"00000E9C";
      when 5904 => data_o <= x"FF005C10";
      when 5905 => data_o <= x"756F74C7";
      when 5906 => data_o <= x"72657070";
      when 5907 => data_o <= x"08FF000C";
      when 5908 => data_o <= x"090012AC";
      when 5909 => data_o <= x"00000EB0";
      when 5910 => data_o <= x"FF005C40";
      when 5911 => data_o <= x"676964C6";
      when 5912 => data_o <= x"FF3F7469";
      when 5913 => data_o <= x"08FF000F";
      when 5914 => data_o <= x"100012AC";
      when 5915 => data_o <= x"00000EE0";
      when 5916 => data_o <= x"FF005C58";
      when 5917 => data_o <= x"756E3EC7";
      when 5918 => data_o <= x"7265626D";
      when 5919 => data_o <= x"08FF0002";
      when 5920 => data_o <= x"170012AC";
      when 5921 => data_o <= x"00000F1C";
      when 5922 => data_o <= x"FF005C70";
      when 5923 => data_o <= x"756F73C6";
      when 5924 => data_o <= x"FF656372";
      when 5925 => data_o <= x"08FF0003";
      when 5926 => data_o <= x"180012AC";
      when 5927 => data_o <= x"00000F24";
      when 5928 => data_o <= x"FF005C88";
      when 5929 => data_o <= x"6F732FC7";
      when 5930 => data_o <= x"65637275";
      when 5931 => data_o <= x"08FF0008";
      when 5932 => data_o <= x"1A0012AC";
      when 5933 => data_o <= x"00000F30";
      when 5934 => data_o <= x"FF005CA0";
      when 5935 => data_o <= x"696B73C4";
      when 5936 => data_o <= x"FFFFFF70";
      when 5937 => data_o <= x"08FF0008";
      when 5938 => data_o <= x"220012AC";
      when 5939 => data_o <= x"00000F50";
      when 5940 => data_o <= x"FF005CB8";
      when 5941 => data_o <= x"616373C4";
      when 5942 => data_o <= x"FFFFFF6E";
      when 5943 => data_o <= x"08FF000A";
      when 5944 => data_o <= x"2A0012AC";
      when 5945 => data_o <= x"00000F70";
      when 5946 => data_o <= x"FF005CD0";
      when 5947 => data_o <= x"726170C5";
      when 5948 => data_o <= x"FFFF6573";
      when 5949 => data_o <= x"08FF0007";
      when 5950 => data_o <= x"2F0012AC";
      when 5951 => data_o <= x"00000F98";
      when 5952 => data_o <= x"FF005CE8";
      when 5953 => data_o <= x"61705FC6";
      when 5954 => data_o <= x"FF657372";
      when 5955 => data_o <= x"08FF0002";
      when 5956 => data_o <= x"330012AC";
      when 5957 => data_o <= x"00000FB4";
      when 5958 => data_o <= x"FF005D00";
      when 5959 => data_o <= x"726170CA";
      when 5960 => data_o <= x"6E2D6573";
      when 5961 => data_o <= x"FF656D61";
      when 5962 => data_o <= x"08FF0005";
      when 5963 => data_o <= x"360012AC";
      when 5964 => data_o <= x"00000FBC";
      when 5965 => data_o <= x"FF005D18";
      when 5966 => data_o <= x"726F77C4";
      when 5967 => data_o <= x"FFFFFF64";
      when 5968 => data_o <= x"08FF0003";
      when 5969 => data_o <= x"3B0012AC";
      when 5970 => data_o <= x"00000FD0";
      when 5971 => data_o <= x"FF005D34";
      when 5972 => data_o <= x"FF282EC2";
      when 5973 => data_o <= x"08FF0002";
      when 5974 => data_o <= x"3E0012AC";
      when 5975 => data_o <= x"00000FDC";
      when 5976 => data_o <= x"FF005D4C";
      when 5977 => data_o <= x"616863C4";
      when 5978 => data_o <= x"FFFFFF72";
      when 5979 => data_o <= x"08FF0012";
      when 5980 => data_o <= x"480012AC";
      when 5981 => data_o <= x"00000FE4";
      when 5982 => data_o <= x"FF005D60";
      when 5983 => data_o <= x"74616DC5";
      when 5984 => data_o <= x"FFFF6863";
      when 5985 => data_o <= x"08FF000E";
      when 5986 => data_o <= x"580012AC";
      when 5987 => data_o <= x"0000102C";
      when 5988 => data_o <= x"FF005D78";
      when 5989 => data_o <= x"66685FC6";
      when 5990 => data_o <= x"FF646E69";
      when 5991 => data_o <= x"08FF000D";
      when 5992 => data_o <= x"630012AC";
      when 5993 => data_o <= x"00001064";
      when 5994 => data_o <= x"FF005D90";
      when 5995 => data_o <= x"696668C5";
      when 5996 => data_o <= x"FFFF646E";
      when 5997 => data_o <= x"08FF0003";
      when 5998 => data_o <= x"6E0012AC";
      when 5999 => data_o <= x"00001098";
      when 6000 => data_o <= x"FF005DA8";
      when 6001 => data_o <= x"736143CF";
      when 6002 => data_o <= x"736E4965";
      when 6003 => data_o <= x"69736E65";
      when 6004 => data_o <= x"65766974";
      when 6005 => data_o <= x"08FF0003";
      when 6006 => data_o <= x"6F0012AC";
      when 6007 => data_o <= x"000010A4";
      when 6008 => data_o <= x"FF005DC0";
      when 6009 => data_o <= x"736143CD";
      when 6010 => data_o <= x"6E655365";
      when 6011 => data_o <= x"69746973";
      when 6012 => data_o <= x"FFFF6576";
      when 6013 => data_o <= x"08FF0004";
      when 6014 => data_o <= x"740012AC";
      when 6015 => data_o <= x"000010B0";
      when 6016 => data_o <= x"FF005DE0";
      when 6017 => data_o <= x"FF2768C2";
      when 6018 => data_o <= x"08FF0002";
      when 6019 => data_o <= x"780012AC";
      when 6020 => data_o <= x"000010C0";
      when 6021 => data_o <= x"FF005E00";
      when 6022 => data_o <= x"FFFF27C1";
      when 6023 => data_o <= x"08FF0006";
      when 6024 => data_o <= x"860012AC";
      when 6025 => data_o <= x"000010C8";
      when 6026 => data_o <= x"FF005E14";
      when 6027 => data_o <= x"6D756ECA";
      when 6028 => data_o <= x"73726562";
      when 6029 => data_o <= x"FF6E6769";
      when 6030 => data_o <= x"08FF0006";
      when 6031 => data_o <= x"8B0012AC";
      when 6032 => data_o <= x"000010E0";
      when 6033 => data_o <= x"FF005E28";
      when 6034 => data_o <= x"6E6F74C8";
      when 6035 => data_o <= x"65626D75";
      when 6036 => data_o <= x"FFFFFF72";
      when 6037 => data_o <= x"08FF0008";
      when 6038 => data_o <= x"900012AC";
      when 6039 => data_o <= x"000010F8";
      when 6040 => data_o <= x"FF005E44";
      when 6041 => data_o <= x"78656EC8";
      when 6042 => data_o <= x"66747574";
      when 6043 => data_o <= x"FFFFFF38";
      when 6044 => data_o <= x"08FF0019";
      when 6045 => data_o <= x"950012AC";
      when 6046 => data_o <= x"00001118";
      when 6047 => data_o <= x"FF005E60";
      when 6048 => data_o <= x"757369C6";
      when 6049 => data_o <= x"FF386674";
      when 6050 => data_o <= x"08FF0028";
      when 6051 => data_o <= x"A50012AC";
      when 6052 => data_o <= x"0000117C";
      when 6053 => data_o <= x"FF005E7C";
      when 6054 => data_o <= x"6E7369C8";
      when 6055 => data_o <= x"65626D75";
      when 6056 => data_o <= x"FFFFFF72";
      when 6057 => data_o <= x"08FF001C";
      when 6058 => data_o <= x"BB0012AC";
      when 6059 => data_o <= x"0000121C";
      when 6060 => data_o <= x"FF005E94";
      when 6061 => data_o <= x"746E69C9";
      when 6062 => data_o <= x"72707265";
      when 6063 => data_o <= x"FFFF7465";
      when 6064 => data_o <= x"00005FB0";
      when 6065 => data_o <= x"2F2E2E12";
      when 6066 => data_o <= x"662F2E2E";
      when 6067 => data_o <= x"6874726F";
      when 6068 => data_o <= x"6165772F";
      when 6069 => data_o <= x"FF662E6E";
      when 6070 => data_o <= x"09FF0003";
      when 6071 => data_o <= x"050012AC";
      when 6072 => data_o <= x"0000128C";
      when 6073 => data_o <= x"FF005EB0";
      when 6074 => data_o <= x"746567C7";
      when 6075 => data_o <= x"6574782D";
      when 6076 => data_o <= x"09FF0001";
      when 6077 => data_o <= x"0F0012AC";
      when 6078 => data_o <= x"000012A4";
      when 6079 => data_o <= x"FF005EE4";
      when 6080 => data_o <= x"2D6F64CC";
      when 6081 => data_o <= x"656D6D69";
      when 6082 => data_o <= x"74616964";
      when 6083 => data_o <= x"FFFFFF65";
      when 6084 => data_o <= x"09FF0001";
      when 6085 => data_o <= x"100012AC";
      when 6086 => data_o <= x"000012A8";
      when 6087 => data_o <= x"FF005EFC";
      when 6088 => data_o <= x"746567C9";
      when 6089 => data_o <= x"63616D2D";
      when 6090 => data_o <= x"FFFF6F72";
      when 6091 => data_o <= x"09FF0001";
      when 6092 => data_o <= x"110012AC";
      when 6093 => data_o <= x"000012AC";
      when 6094 => data_o <= x"FF005F1C";
      when 6095 => data_o <= x"746567CB";
      when 6096 => data_o <= x"6D6F632D";
      when 6097 => data_o <= x"656C6970";
      when 6098 => data_o <= x"09FF0001";
      when 6099 => data_o <= x"120012AC";
      when 6100 => data_o <= x"000012B0";
      when 6101 => data_o <= x"FF005F38";
      when 6102 => data_o <= x"2D6F64C9";
      when 6103 => data_o <= x"73656F64";
      when 6104 => data_o <= x"FFFF652D";
      when 6105 => data_o <= x"09FF0001";
      when 6106 => data_o <= x"130012AC";
      when 6107 => data_o <= x"000012B4";
      when 6108 => data_o <= x"FF005F54";
      when 6109 => data_o <= x"2D6F64C9";
      when 6110 => data_o <= x"73656F64";
      when 6111 => data_o <= x"FFFF632D";
      when 6112 => data_o <= x"09FF0001";
      when 6113 => data_o <= x"140012AC";
      when 6114 => data_o <= x"000012B8";
      when 6115 => data_o <= x"FF005F70";
      when 6116 => data_o <= x"757165C6";
      when 6117 => data_o <= x"FF65655F";
      when 6118 => data_o <= x"09FF0001";
      when 6119 => data_o <= x"150012AC";
      when 6120 => data_o <= x"000012BC";
      when 6121 => data_o <= x"FF005F8C";
      when 6122 => data_o <= x"757165C6";
      when 6123 => data_o <= x"FF63655F";
      when 6124 => data_o <= x"00006240";
      when 6125 => data_o <= x"2F2E2E14";
      when 6126 => data_o <= x"662F2E2E";
      when 6127 => data_o <= x"6874726F";
      when 6128 => data_o <= x"6665642F";
      when 6129 => data_o <= x"2E656E69";
      when 6130 => data_o <= x"FFFFFF66";
      when 6131 => data_o <= x"0AFF0004";
      when 6132 => data_o <= x"030012AC";
      when 6133 => data_o <= x"00001484";
      when 6134 => data_o <= x"FF005FA4";
      when 6135 => data_o <= x"696C61C6";
      when 6136 => data_o <= x"FF686E67";
      when 6137 => data_o <= x"0AFF0004";
      when 6138 => data_o <= x"040012AC";
      when 6139 => data_o <= x"00001494";
      when 6140 => data_o <= x"FF005FD8";
      when 6141 => data_o <= x"696C61C6";
      when 6142 => data_o <= x"FF636E67";
      when 6143 => data_o <= x"0AFF0004";
      when 6144 => data_o <= x"050012AC";
      when 6145 => data_o <= x"000014A4";
      when 6146 => data_o <= x"FF005FF0";
      when 6147 => data_o <= x"696C61C5";
      when 6148 => data_o <= x"FFFF6E67";
      when 6149 => data_o <= x"0AFF0014";
      when 6150 => data_o <= x"140012AC";
      when 6151 => data_o <= x"000014B4";
      when 6152 => data_o <= x"FF006008";
      when 6153 => data_o <= x"616568C7";
      when 6154 => data_o <= x"5B726564";
      when 6155 => data_o <= x"0AFF000E";
      when 6156 => data_o <= x"1F0012AC";
      when 6157 => data_o <= x"00001504";
      when 6158 => data_o <= x"FF006020";
      when 6159 => data_o <= x"65685DC7";
      when 6160 => data_o <= x"72656461";
      when 6161 => data_o <= x"0AFF0002";
      when 6162 => data_o <= x"260012AC";
      when 6163 => data_o <= x"0000153C";
      when 6164 => data_o <= x"FF006038";
      when 6165 => data_o <= x"616C66C6";
      when 6166 => data_o <= x"FF217367";
      when 6167 => data_o <= x"0AFF0005";
      when 6168 => data_o <= x"310012AC";
      when 6169 => data_o <= x"00001544";
      when 6170 => data_o <= x"FF006050";
      when 6171 => data_o <= x"757165C3";
      when 6172 => data_o <= x"0AFF0002";
      when 6173 => data_o <= x"370012AC";
      when 6174 => data_o <= x"00001558";
      when 6175 => data_o <= x"FF006068";
      when 6176 => data_o <= x"73616CC4";
      when 6177 => data_o <= x"FFFFFF74";
      when 6178 => data_o <= x"0AFF0002";
      when 6179 => data_o <= x"380012AC";
      when 6180 => data_o <= x"00001560";
      when 6181 => data_o <= x"FF00607C";
      when 6182 => data_o <= x"726C63C7";
      when 6183 => data_o <= x"7473616C";
      when 6184 => data_o <= x"0AFF0002";
      when 6185 => data_o <= x"390012AC";
      when 6186 => data_o <= x"00001568";
      when 6187 => data_o <= x"FF006094";
      when 6188 => data_o <= x"726C63CB";
      when 6189 => data_o <= x"6374782D";
      when 6190 => data_o <= x"73746962";
      when 6191 => data_o <= x"0AFF0002";
      when 6192 => data_o <= x"3B0012AC";
      when 6193 => data_o <= x"00001570";
      when 6194 => data_o <= x"FF0060AC";
      when 6195 => data_o <= x"726C63CC";
      when 6196 => data_o <= x"616C662D";
      when 6197 => data_o <= x"74696267";
      when 6198 => data_o <= x"FFFFFF73";
      when 6199 => data_o <= x"0AFF0002";
      when 6200 => data_o <= x"3C0012AC";
      when 6201 => data_o <= x"00001578";
      when 6202 => data_o <= x"FF0060C8";
      when 6203 => data_o <= x"63616DC5";
      when 6204 => data_o <= x"FFFF6F72";
      when 6205 => data_o <= x"0AFF0002";
      when 6206 => data_o <= x"3D0012AC";
      when 6207 => data_o <= x"00001580";
      when 6208 => data_o <= x"FF0060E8";
      when 6209 => data_o <= x"6D6D69C9";
      when 6210 => data_o <= x"61696465";
      when 6211 => data_o <= x"FFFF6574";
      when 6212 => data_o <= x"0AFF0002";
      when 6213 => data_o <= x"3E0012AC";
      when 6214 => data_o <= x"00001588";
      when 6215 => data_o <= x"FF006100";
      when 6216 => data_o <= x"6C6163C9";
      when 6217 => data_o <= x"6E6F2D6C";
      when 6218 => data_o <= x"FFFF796C";
      when 6219 => data_o <= x"0AFF0003";
      when 6220 => data_o <= x"400012AC";
      when 6221 => data_o <= x"00001590";
      when 6222 => data_o <= x"FF00611C";
      when 6223 => data_o <= x"FFFF5DC1";
      when 6224 => data_o <= x"0AFF0003";
      when 6225 => data_o <= x"410012A4";
      when 6226 => data_o <= x"0000159C";
      when 6227 => data_o <= x"FF006138";
      when 6228 => data_o <= x"FFFF5BC1";
      when 6229 => data_o <= x"0AFF0019";
      when 6230 => data_o <= x"430012A4";
      when 6231 => data_o <= x"000015A8";
      when 6232 => data_o <= x"FF00614C";
      when 6233 => data_o <= x"FFFF3BC1";
      when 6234 => data_o <= x"0AFF000B";
      when 6235 => data_o <= x"500012AC";
      when 6236 => data_o <= x"0000160C";
      when 6237 => data_o <= x"FF006160";
      when 6238 => data_o <= x"FF3A2BC2";
      when 6239 => data_o <= x"0AFF0002";
      when 6240 => data_o <= x"580012AC";
      when 6241 => data_o <= x"00001638";
      when 6242 => data_o <= x"FF006174";
      when 6243 => data_o <= x"FFFF3AC1";
      when 6244 => data_o <= x"0AFF0004";
      when 6245 => data_o <= x"5B0012AC";
      when 6246 => data_o <= x"00001640";
      when 6247 => data_o <= x"00006188";
      when 6248 => data_o <= x"6F6E3AC7";
      when 6249 => data_o <= x"656D616E";
      when 6250 => data_o <= x"0AFF0002";
      when 6251 => data_o <= x"6A0012AC";
      when 6252 => data_o <= x"00001650";
      when 6253 => data_o <= x"0000619C";
      when 6254 => data_o <= x"726568C4";
      when 6255 => data_o <= x"FFFFFF65";
      when 6256 => data_o <= x"0AFF0002";
      when 6257 => data_o <= x"6B0012AC";
      when 6258 => data_o <= x"00001658";
      when 6259 => data_o <= x"000061B4";
      when 6260 => data_o <= x"6C6C61C5";
      when 6261 => data_o <= x"FFFF746F";
      when 6262 => data_o <= x"0AFF0004";
      when 6263 => data_o <= x"6C0012AC";
      when 6264 => data_o <= x"00001660";
      when 6265 => data_o <= x"000061CC";
      when 6266 => data_o <= x"6C612FC6";
      when 6267 => data_o <= x"FF746F6C";
      when 6268 => data_o <= x"0AFF0003";
      when 6269 => data_o <= x"6D0012AC";
      when 6270 => data_o <= x"00001670";
      when 6271 => data_o <= x"000061E4";
      when 6272 => data_o <= x"667562C7";
      when 6273 => data_o <= x"3A726566";
      when 6274 => data_o <= x"0AFF0001";
      when 6275 => data_o <= x"6E0012AC";
      when 6276 => data_o <= x"0000167C";
      when 6277 => data_o <= x"000061FC";
      when 6278 => data_o <= x"6E6F63C8";
      when 6279 => data_o <= x"6E617473";
      when 6280 => data_o <= x"FFFFFF74";
      when 6281 => data_o <= x"0AFF0005";
      when 6282 => data_o <= x"6F0012AC";
      when 6283 => data_o <= x"00001680";
      when 6284 => data_o <= x"00006214";
      when 6285 => data_o <= x"726176C8";
      when 6286 => data_o <= x"6C626169";
      when 6287 => data_o <= x"FFFFFF65";
      when 6288 => data_o <= x"000067EC";
      when 6289 => data_o <= x"2F2E2E17";
      when 6290 => data_o <= x"662F2E2E";
      when 6291 => data_o <= x"6874726F";
      when 6292 => data_o <= x"7274732F";
      when 6293 => data_o <= x"75746375";
      when 6294 => data_o <= x"662E6572";
      when 6295 => data_o <= x"0BFF0003";
      when 6296 => data_o <= x"030012A4";
      when 6297 => data_o <= x"00001694";
      when 6298 => data_o <= x"00006230";
      when 6299 => data_o <= x"FFFF5CC1";
      when 6300 => data_o <= x"0BFF0001";
      when 6301 => data_o <= x"040012A4";
      when 6302 => data_o <= x"000016A0";
      when 6303 => data_o <= x"00006268";
      when 6304 => data_o <= x"74696CC7";
      when 6305 => data_o <= x"6C617265";
      when 6306 => data_o <= x"0BFF0002";
      when 6307 => data_o <= x"050012A4";
      when 6308 => data_o <= x"000016A4";
      when 6309 => data_o <= x"0000627C";
      when 6310 => data_o <= x"68635BC6";
      when 6311 => data_o <= x"FF5D7261";
      when 6312 => data_o <= x"0BFF0001";
      when 6313 => data_o <= x"060012A4";
      when 6314 => data_o <= x"000016AC";
      when 6315 => data_o <= x"00006294";
      when 6316 => data_o <= x"697865C4";
      when 6317 => data_o <= x"FFFFFF74";
      when 6318 => data_o <= x"0BFF0001";
      when 6319 => data_o <= x"070012A4";
      when 6320 => data_o <= x"000016B0";
      when 6321 => data_o <= x"000062AC";
      when 6322 => data_o <= x"616863C5";
      when 6323 => data_o <= x"FFFF7372";
      when 6324 => data_o <= x"0BFF0003";
      when 6325 => data_o <= x"080012A4";
      when 6326 => data_o <= x"000016B4";
      when 6327 => data_o <= x"000062C4";
      when 6328 => data_o <= x"FFFF28C1";
      when 6329 => data_o <= x"0BFF0002";
      when 6330 => data_o <= x"0B0012A4";
      when 6331 => data_o <= x"000016C0";
      when 6332 => data_o <= x"000062DC";
      when 6333 => data_o <= x"5D275BC3";
      when 6334 => data_o <= x"0BFF0004";
      when 6335 => data_o <= x"0F0012AC";
      when 6336 => data_o <= x"000016C8";
      when 6337 => data_o <= x"000062F0";
      when 6338 => data_o <= x"657478C6";
      when 6339 => data_o <= x"FF637478";
      when 6340 => data_o <= x"0BFF0003";
      when 6341 => data_o <= x"120012AC";
      when 6342 => data_o <= x"000016D8";
      when 6343 => data_o <= x"00006304";
      when 6344 => data_o <= x"667478C6";
      when 6345 => data_o <= x"FF67616C";
      when 6346 => data_o <= x"0BFF0004";
      when 6347 => data_o <= x"150012AC";
      when 6348 => data_o <= x"000016E4";
      when 6349 => data_o <= x"0000631C";
      when 6350 => data_o <= x"616573CF";
      when 6351 => data_o <= x"2D686372";
      when 6352 => data_o <= x"64726F77";
      when 6353 => data_o <= x"7473696C";
      when 6354 => data_o <= x"0BFF0009";
      when 6355 => data_o <= x"1A0012A4";
      when 6356 => data_o <= x"000016F4";
      when 6357 => data_o <= x"00006334";
      when 6358 => data_o <= x"736F70C8";
      when 6359 => data_o <= x"6E6F7074";
      when 6360 => data_o <= x"FFFFFF65";
      when 6361 => data_o <= x"0BFF0004";
      when 6362 => data_o <= x"210012A4";
      when 6363 => data_o <= x"00001718";
      when 6364 => data_o <= x"00006354";
      when 6365 => data_o <= x"636572C7";
      when 6366 => data_o <= x"65737275";
      when 6367 => data_o <= x"0BFF0003";
      when 6368 => data_o <= x"290012AC";
      when 6369 => data_o <= x"00001728";
      when 6370 => data_o <= x"00006370";
      when 6371 => data_o <= x"456F4EC9";
      when 6372 => data_o <= x"75636578";
      when 6373 => data_o <= x"FFFF6574";
      when 6374 => data_o <= x"0BFF000D";
      when 6375 => data_o <= x"2C0012AC";
      when 6376 => data_o <= x"00001734";
      when 6377 => data_o <= x"00006388";
      when 6378 => data_o <= x"65654EC8";
      when 6379 => data_o <= x"6F6C5364";
      when 6380 => data_o <= x"FFFFFF74";
      when 6381 => data_o <= x"0BFF0002";
      when 6382 => data_o <= x"330012AC";
      when 6383 => data_o <= x"00001768";
      when 6384 => data_o <= x"000063A4";
      when 6385 => data_o <= x"72625FC7";
      when 6386 => data_o <= x"68636E61";
      when 6387 => data_o <= x"0BFF0009";
      when 6388 => data_o <= x"360012AC";
      when 6389 => data_o <= x"00001770";
      when 6390 => data_o <= x"000063C0";
      when 6391 => data_o <= x"756A5FC5";
      when 6392 => data_o <= x"FFFF706D";
      when 6393 => data_o <= x"0BFF0011";
      when 6394 => data_o <= x"3B0012A4";
      when 6395 => data_o <= x"00001794";
      when 6396 => data_o <= x"000063D8";
      when 6397 => data_o <= x"656874C4";
      when 6398 => data_o <= x"FFFFFF6E";
      when 6399 => data_o <= x"0BFF0006";
      when 6400 => data_o <= x"450012A4";
      when 6401 => data_o <= x"000017D8";
      when 6402 => data_o <= x"000063F0";
      when 6403 => data_o <= x"676562C5";
      when 6404 => data_o <= x"FFFF6E69";
      when 6405 => data_o <= x"0BFF0009";
      when 6406 => data_o <= x"4A0012A4";
      when 6407 => data_o <= x"000017F0";
      when 6408 => data_o <= x"00006408";
      when 6409 => data_o <= x"616761C5";
      when 6410 => data_o <= x"FFFF6E69";
      when 6411 => data_o <= x"0BFF0003";
      when 6412 => data_o <= x"530012A4";
      when 6413 => data_o <= x"00001814";
      when 6414 => data_o <= x"00006420";
      when 6415 => data_o <= x"656861C5";
      when 6416 => data_o <= x"FFFF6461";
      when 6417 => data_o <= x"0BFF0005";
      when 6418 => data_o <= x"560012A4";
      when 6419 => data_o <= x"00001820";
      when 6420 => data_o <= x"00006438";
      when 6421 => data_o <= x"6E6669C4";
      when 6422 => data_o <= x"FFFFFF63";
      when 6423 => data_o <= x"0BFF0005";
      when 6424 => data_o <= x"5A0012A4";
      when 6425 => data_o <= x"00001834";
      when 6426 => data_o <= x"00006450";
      when 6427 => data_o <= x"FF6669C2";
      when 6428 => data_o <= x"0BFF0005";
      when 6429 => data_o <= x"5E0012A4";
      when 6430 => data_o <= x"00001848";
      when 6431 => data_o <= x"00006468";
      when 6432 => data_o <= x"66692BC3";
      when 6433 => data_o <= x"0BFF0002";
      when 6434 => data_o <= x"620012A4";
      when 6435 => data_o <= x"0000185C";
      when 6436 => data_o <= x"0000647C";
      when 6437 => data_o <= x"736C65C4";
      when 6438 => data_o <= x"FFFFFF65";
      when 6439 => data_o <= x"0BFF0003";
      when 6440 => data_o <= x"660012A4";
      when 6441 => data_o <= x"00001864";
      when 6442 => data_o <= x"00006490";
      when 6443 => data_o <= x"696877C5";
      when 6444 => data_o <= x"FFFF656C";
      when 6445 => data_o <= x"0BFF0003";
      when 6446 => data_o <= x"690012A4";
      when 6447 => data_o <= x"00001870";
      when 6448 => data_o <= x"000064A8";
      when 6449 => data_o <= x"68772BC6";
      when 6450 => data_o <= x"FF656C69";
      when 6451 => data_o <= x"0BFF0002";
      when 6452 => data_o <= x"6C0012A4";
      when 6453 => data_o <= x"0000187C";
      when 6454 => data_o <= x"000064C0";
      when 6455 => data_o <= x"706572C6";
      when 6456 => data_o <= x"FF746165";
      when 6457 => data_o <= x"0BFF0005";
      when 6458 => data_o <= x"700012A4";
      when 6459 => data_o <= x"00001884";
      when 6460 => data_o <= x"000064D8";
      when 6461 => data_o <= x"6E752BC6";
      when 6462 => data_o <= x"FF6C6974";
      when 6463 => data_o <= x"0BFF0005";
      when 6464 => data_o <= x"750012A4";
      when 6465 => data_o <= x"00001898";
      when 6466 => data_o <= x"000064F0";
      when 6467 => data_o <= x"746E75C5";
      when 6468 => data_o <= x"FFFF6C69";
      when 6469 => data_o <= x"0BFF0004";
      when 6470 => data_o <= x"7A0012A4";
      when 6471 => data_o <= x"000018AC";
      when 6472 => data_o <= x"00006508";
      when 6473 => data_o <= x"6F6672C4";
      when 6474 => data_o <= x"FFFFFF72";
      when 6475 => data_o <= x"0BFF0003";
      when 6476 => data_o <= x"7E0012A4";
      when 6477 => data_o <= x"000018BC";
      when 6478 => data_o <= x"00006520";
      when 6479 => data_o <= x"726F66C3";
      when 6480 => data_o <= x"0BFF0002";
      when 6481 => data_o <= x"820012A4";
      when 6482 => data_o <= x"000018C8";
      when 6483 => data_o <= x"00006538";
      when 6484 => data_o <= x"78656EC4";
      when 6485 => data_o <= x"FFFFFF74";
      when 6486 => data_o <= x"0BFF0009";
      when 6487 => data_o <= x"890012AC";
      when 6488 => data_o <= x"000018D0";
      when 6489 => data_o <= x"0000654C";
      when 6490 => data_o <= x"72635FC7";
      when 6491 => data_o <= x"65746165";
      when 6492 => data_o <= x"0BFF0006";
      when 6493 => data_o <= x"8F0012AC";
      when 6494 => data_o <= x"000018F4";
      when 6495 => data_o <= x"00006564";
      when 6496 => data_o <= x"666564C5";
      when 6497 => data_o <= x"FFFF7265";
      when 6498 => data_o <= x"0BFF0005";
      when 6499 => data_o <= x"930012AC";
      when 6500 => data_o <= x"0000190C";
      when 6501 => data_o <= x"0000657C";
      when 6502 => data_o <= x"FF7369C2";
      when 6503 => data_o <= x"0BFF0010";
      when 6504 => data_o <= x"960012AC";
      when 6505 => data_o <= x"00001920";
      when 6506 => data_o <= x"00006594";
      when 6507 => data_o <= x"657263C6";
      when 6508 => data_o <= x"FF657461";
      when 6509 => data_o <= x"0BFF0005";
      when 6510 => data_o <= x"9F0012AC";
      when 6511 => data_o <= x"00001960";
      when 6512 => data_o <= x"000065A8";
      when 6513 => data_o <= x"637369C6";
      when 6514 => data_o <= x"FF3F6D6F";
      when 6515 => data_o <= x"0BFF0009";
      when 6516 => data_o <= x"A40012AC";
      when 6517 => data_o <= x"00001974";
      when 6518 => data_o <= x"000065C0";
      when 6519 => data_o <= x"623E5FC6";
      when 6520 => data_o <= x"FF79646F";
      when 6521 => data_o <= x"0BFF0002";
      when 6522 => data_o <= x"AE0012AC";
      when 6523 => data_o <= x"00001998";
      when 6524 => data_o <= x"000065D8";
      when 6525 => data_o <= x"6F623EC5";
      when 6526 => data_o <= x"FFFF7964";
      when 6527 => data_o <= x"0BFF000C";
      when 6528 => data_o <= x"B70012AC";
      when 6529 => data_o <= x"000019A0";
      when 6530 => data_o <= x"000065F0";
      when 6531 => data_o <= x"656F64C5";
      when 6532 => data_o <= x"FFFF3E73";
      when 6533 => data_o <= x"0BFF0002";
      when 6534 => data_o <= x"C60012A4";
      when 6535 => data_o <= x"000019D0";
      when 6536 => data_o <= x"00006608";
      when 6537 => data_o <= x"736163C4";
      when 6538 => data_o <= x"FFFFFF65";
      when 6539 => data_o <= x"0BFF0003";
      when 6540 => data_o <= x"C90012A4";
      when 6541 => data_o <= x"000019D8";
      when 6542 => data_o <= x"00006620";
      when 6543 => data_o <= x"FF666FC2";
      when 6544 => data_o <= x"0BFF0001";
      when 6545 => data_o <= x"CC0012A4";
      when 6546 => data_o <= x"000019E4";
      when 6547 => data_o <= x"00006638";
      when 6548 => data_o <= x"646E65C5";
      when 6549 => data_o <= x"FFFF666F";
      when 6550 => data_o <= x"0BFF0007";
      when 6551 => data_o <= x"CF0012A4";
      when 6552 => data_o <= x"000019E8";
      when 6553 => data_o <= x"0000664C";
      when 6554 => data_o <= x"646E65C7";
      when 6555 => data_o <= x"65736163";
      when 6556 => data_o <= x"0BFF0010";
      when 6557 => data_o <= x"D80012A4";
      when 6558 => data_o <= x"00001A04";
      when 6559 => data_o <= x"00006664";
      when 6560 => data_o <= x"FF6F64C2";
      when 6561 => data_o <= x"0BFF0008";
      when 6562 => data_o <= x"DE0012A4";
      when 6563 => data_o <= x"00001A44";
      when 6564 => data_o <= x"0000667C";
      when 6565 => data_o <= x"6F643FC3";
      when 6566 => data_o <= x"0BFF0004";
      when 6567 => data_o <= x"E40012AC";
      when 6568 => data_o <= x"00001A64";
      when 6569 => data_o <= x"00006690";
      when 6570 => data_o <= x"737570C6";
      when 6571 => data_o <= x"FF564C68";
      when 6572 => data_o <= x"0BFF0005";
      when 6573 => data_o <= x"E50012AC";
      when 6574 => data_o <= x"00001A74";
      when 6575 => data_o <= x"000066A4";
      when 6576 => data_o <= x"706F70C5";
      when 6577 => data_o <= x"FFFF564C";
      when 6578 => data_o <= x"0BFF0005";
      when 6579 => data_o <= x"E70012A4";
      when 6580 => data_o <= x"00001A88";
      when 6581 => data_o <= x"000066BC";
      when 6582 => data_o <= x"61656CC5";
      when 6583 => data_o <= x"FFFF6576";
      when 6584 => data_o <= x"0BFF0007";
      when 6585 => data_o <= x"EB0012AC";
      when 6586 => data_o <= x"00001A9C";
      when 6587 => data_o <= x"000066D4";
      when 6588 => data_o <= x"656C5FC7";
      when 6589 => data_o <= x"73657661";
      when 6590 => data_o <= x"0BFF0005";
      when 6591 => data_o <= x"F00012A4";
      when 6592 => data_o <= x"00001AB8";
      when 6593 => data_o <= x"000066EC";
      when 6594 => data_o <= x"6F6F6CC4";
      when 6595 => data_o <= x"FFFFFF70";
      when 6596 => data_o <= x"0BFF0005";
      when 6597 => data_o <= x"F30012A4";
      when 6598 => data_o <= x"00001ACC";
      when 6599 => data_o <= x"00006704";
      when 6600 => data_o <= x"6F6C2BC5";
      when 6601 => data_o <= x"FFFF706F";
      when 6602 => data_o <= x"0BFF0003";
      when 6603 => data_o <= x"F60012A4";
      when 6604 => data_o <= x"00001AE0";
      when 6605 => data_o <= x"0000671C";
      when 6606 => data_o <= x"FFFF69C1";
      when 6607 => data_o <= x"0BFF0008";
      when 6608 => data_o <= x"FC0012AC";
      when 6609 => data_o <= x"00001AEC";
      when 6610 => data_o <= x"00006734";
      when 6611 => data_o <= x"FF222CC2";
      when 6612 => data_o <= x"0BFF0004";
      when 6613 => data_o <= x"020012AC";
      when 6614 => data_o <= x"01001B0C";
      when 6615 => data_o <= x"00006748";
      when 6616 => data_o <= x"22785FC3";
      when 6617 => data_o <= x"0BFF0005";
      when 6618 => data_o <= x"050012A4";
      when 6619 => data_o <= x"01001B1C";
      when 6620 => data_o <= x"0000675C";
      when 6621 => data_o <= x"FF222EC2";
      when 6622 => data_o <= x"0BFF0002";
      when 6623 => data_o <= x"0A0012AC";
      when 6624 => data_o <= x"01001B30";
      when 6625 => data_o <= x"00006770";
      when 6626 => data_o <= x"6F6261C5";
      when 6627 => data_o <= x"FFFF7472";
      when 6628 => data_o <= x"0BFF0005";
      when 6629 => data_o <= x"0C0012A4";
      when 6630 => data_o <= x"01001B38";
      when 6631 => data_o <= x"00006784";
      when 6632 => data_o <= x"6F6261C6";
      when 6633 => data_o <= x"FF227472";
      when 6634 => data_o <= x"0BFF0007";
      when 6635 => data_o <= x"170012AC";
      when 6636 => data_o <= x"01001B4C";
      when 6637 => data_o <= x"0000679C";
      when 6638 => data_o <= x"617274CA";
      when 6639 => data_o <= x"6569736E";
      when 6640 => data_o <= x"FF22746E";
      when 6641 => data_o <= x"0BFF0002";
      when 6642 => data_o <= x"20001B68";
      when 6643 => data_o <= x"01001B74";
      when 6644 => data_o <= x"000067B4";
      when 6645 => data_o <= x"FF2253C2";
      when 6646 => data_o <= x"0BFF0001";
      when 6647 => data_o <= x"21001B0C";
      when 6648 => data_o <= x"01001B7C";
      when 6649 => data_o <= x"000067D0";
      when 6650 => data_o <= x"FF2243C2";
      when 6651 => data_o <= x"00006878";
      when 6652 => data_o <= x"2F2E2E16";
      when 6653 => data_o <= x"662F2E2E";
      when 6654 => data_o <= x"6874726F";
      when 6655 => data_o <= x"6176652F";
      when 6656 => data_o <= x"7461756C";
      when 6657 => data_o <= x"FF662E65";
      when 6658 => data_o <= x"0CFF0002";
      when 6659 => data_o <= x"040012AC";
      when 6660 => data_o <= x"00001B80";
      when 6661 => data_o <= x"000067E4";
      when 6662 => data_o <= x"756F73C6";
      when 6663 => data_o <= x"FF656372";
      when 6664 => data_o <= x"0CFF0007";
      when 6665 => data_o <= x"070012AC";
      when 6666 => data_o <= x"00001B88";
      when 6667 => data_o <= x"00006814";
      when 6668 => data_o <= x"766173CA";
      when 6669 => data_o <= x"6E692D65";
      when 6670 => data_o <= x"FF747570";
      when 6671 => data_o <= x"0CFF000D";
      when 6672 => data_o <= x"0C0012AC";
      when 6673 => data_o <= x"00001BA4";
      when 6674 => data_o <= x"0000682C";
      when 6675 => data_o <= x"736572CD";
      when 6676 => data_o <= x"65726F74";
      when 6677 => data_o <= x"706E692D";
      when 6678 => data_o <= x"FFFF7475";
      when 6679 => data_o <= x"0CFF0014";
      when 6680 => data_o <= x"130012AC";
      when 6681 => data_o <= x"00001BD8";
      when 6682 => data_o <= x"00006848";
      when 6683 => data_o <= x"617665C8";
      when 6684 => data_o <= x"7461756C";
      when 6685 => data_o <= x"FFFFFF65";
      when 6686 => data_o <= x"000068F0";
      when 6687 => data_o <= x"2F2E2E12";
      when 6688 => data_o <= x"662F2E2E";
      when 6689 => data_o <= x"6874726F";
      when 6690 => data_o <= x"6975712F";
      when 6691 => data_o <= x"FF662E74";
      when 6692 => data_o <= x"0DFF0014";
      when 6693 => data_o <= x"050012AC";
      when 6694 => data_o <= x"00001C28";
      when 6695 => data_o <= x"00006868";
      when 6696 => data_o <= x"666572C6";
      when 6697 => data_o <= x"FF6C6C69";
      when 6698 => data_o <= x"0DFF0004";
      when 6699 => data_o <= x"0E0012AC";
      when 6700 => data_o <= x"00001C78";
      when 6701 => data_o <= x"0000689C";
      when 6702 => data_o <= x"757128C6";
      when 6703 => data_o <= x"FF297469";
      when 6704 => data_o <= x"0DFF000B";
      when 6705 => data_o <= x"150012AC";
      when 6706 => data_o <= x"00001C88";
      when 6707 => data_o <= x"000068B4";
      when 6708 => data_o <= x"75712EC5";
      when 6709 => data_o <= x"FFFF7469";
      when 6710 => data_o <= x"0DFF0016";
      when 6711 => data_o <= x"1A0012AC";
      when 6712 => data_o <= x"00001CB4";
      when 6713 => data_o <= x"000068CC";
      when 6714 => data_o <= x"697571C4";
      when 6715 => data_o <= x"FFFFFF74";
      when 6716 => data_o <= x"00006B08";
      when 6717 => data_o <= x"2F2E2E13";
      when 6718 => data_o <= x"662F2E2E";
      when 6719 => data_o <= x"6874726F";
      when 6720 => data_o <= x"64726F2F";
      when 6721 => data_o <= x"662E7265";
      when 6722 => data_o <= x"0EFF0016";
      when 6723 => data_o <= x"040012AC";
      when 6724 => data_o <= x"00001D0C";
      when 6725 => data_o <= x"000068E4";
      when 6726 => data_o <= x"6F775FC9";
      when 6727 => data_o <= x"696C6472";
      when 6728 => data_o <= x"FFFF7473";
      when 6729 => data_o <= x"0EFF0002";
      when 6730 => data_o <= x"0F0012AC";
      when 6731 => data_o <= x"00001D64";
      when 6732 => data_o <= x"00006914";
      when 6733 => data_o <= x"726F77C8";
      when 6734 => data_o <= x"73696C64";
      when 6735 => data_o <= x"FFFFFF74";
      when 6736 => data_o <= x"0EFF000A";
      when 6737 => data_o <= x"120012AC";
      when 6738 => data_o <= x"00001D6C";
      when 6739 => data_o <= x"00006930";
      when 6740 => data_o <= x"772E28C6";
      when 6741 => data_o <= x"FF296469";
      when 6742 => data_o <= x"0EFF000D";
      when 6743 => data_o <= x"180012AC";
      when 6744 => data_o <= x"00001D94";
      when 6745 => data_o <= x"0000694C";
      when 6746 => data_o <= x"69772EC4";
      when 6747 => data_o <= x"FFFFFF64";
      when 6748 => data_o <= x"0EFF0006";
      when 6749 => data_o <= x"200012AC";
      when 6750 => data_o <= x"00001DC8";
      when 6751 => data_o <= x"00006964";
      when 6752 => data_o <= x"6E6966C4";
      when 6753 => data_o <= x"FFFFFF64";
      when 6754 => data_o <= x"0EFF000A";
      when 6755 => data_o <= x"260012AC";
      when 6756 => data_o <= x"00001DE0";
      when 6757 => data_o <= x"0000697C";
      when 6758 => data_o <= x"746567C9";
      when 6759 => data_o <= x"64726F2D";
      when 6760 => data_o <= x"FFFF7265";
      when 6761 => data_o <= x"0EFF000E";
      when 6762 => data_o <= x"2B0012AC";
      when 6763 => data_o <= x"00001E08";
      when 6764 => data_o <= x"00006994";
      when 6765 => data_o <= x"746573C9";
      when 6766 => data_o <= x"64726F2D";
      when 6767 => data_o <= x"FFFF7265";
      when 6768 => data_o <= x"0EFF0002";
      when 6769 => data_o <= x"2F0012AC";
      when 6770 => data_o <= x"00001E40";
      when 6771 => data_o <= x"000069B0";
      when 6772 => data_o <= x"746573CB";
      when 6773 => data_o <= x"7275632D";
      when 6774 => data_o <= x"746E6572";
      when 6775 => data_o <= x"0EFF0002";
      when 6776 => data_o <= x"300012AC";
      when 6777 => data_o <= x"00001E48";
      when 6778 => data_o <= x"000069CC";
      when 6779 => data_o <= x"746567CB";
      when 6780 => data_o <= x"7275632D";
      when 6781 => data_o <= x"746E6572";
      when 6782 => data_o <= x"0EFF0002";
      when 6783 => data_o <= x"310012AC";
      when 6784 => data_o <= x"00001E50";
      when 6785 => data_o <= x"000069E8";
      when 6786 => data_o <= x"6C6E6FC4";
      when 6787 => data_o <= x"FFFFFF79";
      when 6788 => data_o <= x"0EFF0003";
      when 6789 => data_o <= x"320012AC";
      when 6790 => data_o <= x"00001E58";
      when 6791 => data_o <= x"00006A04";
      when 6792 => data_o <= x"736C61C4";
      when 6793 => data_o <= x"FFFFFF6F";
      when 6794 => data_o <= x"0EFF0003";
      when 6795 => data_o <= x"340012AC";
      when 6796 => data_o <= x"00001E64";
      when 6797 => data_o <= x"00006A1C";
      when 6798 => data_o <= x"657270C8";
      when 6799 => data_o <= x"756F6976";
      when 6800 => data_o <= x"FFFFFF73";
      when 6801 => data_o <= x"0EFF0003";
      when 6802 => data_o <= x"360012AC";
      when 6803 => data_o <= x"00001E70";
      when 6804 => data_o <= x"00006A34";
      when 6805 => data_o <= x"666564CB";
      when 6806 => data_o <= x"74696E69";
      when 6807 => data_o <= x"736E6F69";
      when 6808 => data_o <= x"0EFF0004";
      when 6809 => data_o <= x"390012AC";
      when 6810 => data_o <= x"00001E7C";
      when 6811 => data_o <= x"00006A50";
      when 6812 => data_o <= x"6F662FC6";
      when 6813 => data_o <= x"FF687472";
      when 6814 => data_o <= x"0EFF0003";
      when 6815 => data_o <= x"3A0012AC";
      when 6816 => data_o <= x"00001E8C";
      when 6817 => data_o <= x"00006A6C";
      when 6818 => data_o <= x"726F66C5";
      when 6819 => data_o <= x"FFFF6874";
      when 6820 => data_o <= x"0EFF0016";
      when 6821 => data_o <= x"3D0012AC";
      when 6822 => data_o <= x"00001E98";
      when 6823 => data_o <= x"00006A84";
      when 6824 => data_o <= x"64726FC5";
      when 6825 => data_o <= x"FFFF7265";
      when 6826 => data_o <= x"0EFF000D";
      when 6827 => data_o <= x"450012AC";
      when 6828 => data_o <= x"00001EF0";
      when 6829 => data_o <= x"00006A9C";
      when 6830 => data_o <= x"657377C7";
      when 6831 => data_o <= x"68637261";
      when 6832 => data_o <= x"0EFF001B";
      when 6833 => data_o <= x"4F0012AC";
      when 6834 => data_o <= x"00001F24";
      when 6835 => data_o <= x"00006AB4";
      when 6836 => data_o <= x"6F775FC6";
      when 6837 => data_o <= x"FF736472";
      when 6838 => data_o <= x"0EFF000B";
      when 6839 => data_o <= x"5D0012AC";
      when 6840 => data_o <= x"00001F90";
      when 6841 => data_o <= x"00006ACC";
      when 6842 => data_o <= x"726F77C5";
      when 6843 => data_o <= x"FFFF7364";
      when 6844 => data_o <= x"0EFF0002";
      when 6845 => data_o <= x"630012AC";
      when 6846 => data_o <= x"00001FBC";
      when 6847 => data_o <= x"00006AE4";
      when 6848 => data_o <= x"6F7777C6";
      when 6849 => data_o <= x"FF736472";
      when 6850 => data_o <= x"00006C78";
      when 6851 => data_o <= x"2F2E2E11";
      when 6852 => data_o <= x"662F2E2E";
      when 6853 => data_o <= x"6874726F";
      when 6854 => data_o <= x"6565732F";
      when 6855 => data_o <= x"FFFF662E";
      when 6856 => data_o <= x"00001FC4";
      when 6857 => data_o <= x"0FFFFFFF";
      when 6858 => data_o <= x"060012BC";
      when 6859 => data_o <= x"000012B8";
      when 6860 => data_o <= x"00006AFC";
      when 6861 => data_o <= x"6E706F07";
      when 6862 => data_o <= x"73656D61";
      when 6863 => data_o <= x"0FFF0006";
      when 6864 => data_o <= x"110012AC";
      when 6865 => data_o <= x"000020A0";
      when 6866 => data_o <= x"00006B30";
      when 6867 => data_o <= x"6E706FC6";
      when 6868 => data_o <= x"FF656D61";
      when 6869 => data_o <= x"000020B8";
      when 6870 => data_o <= x"0FFFFFFF";
      when 6871 => data_o <= x"180012BC";
      when 6872 => data_o <= x"000012B8";
      when 6873 => data_o <= x"00006B48";
      when 6874 => data_o <= x"69706F07";
      when 6875 => data_o <= x"64656D6D";
      when 6876 => data_o <= x"000020C0";
      when 6877 => data_o <= x"0FFFFFFF";
      when 6878 => data_o <= x"1B0012BC";
      when 6879 => data_o <= x"000012B8";
      when 6880 => data_o <= x"00006B64";
      when 6881 => data_o <= x"69706F09";
      when 6882 => data_o <= x"64616D6D";
      when 6883 => data_o <= x"FFFF7264";
      when 6884 => data_o <= x"0FFF000A";
      when 6885 => data_o <= x"210012AC";
      when 6886 => data_o <= x"000020C4";
      when 6887 => data_o <= x"00006B80";
      when 6888 => data_o <= x"697369C5";
      when 6889 => data_o <= x"FFFF6D6D";
      when 6890 => data_o <= x"0FFF0009";
      when 6891 => data_o <= x"2A0012AC";
      when 6892 => data_o <= x"000020EC";
      when 6893 => data_o <= x"00006B9C";
      when 6894 => data_o <= x"74785FC7";
      when 6895 => data_o <= x"656D616E";
      when 6896 => data_o <= x"0FFF000E";
      when 6897 => data_o <= x"320012AC";
      when 6898 => data_o <= x"00002110";
      when 6899 => data_o <= x"00006BB4";
      when 6900 => data_o <= x"6E7478C6";
      when 6901 => data_o <= x"FF656D61";
      when 6902 => data_o <= x"0FFF001D";
      when 6903 => data_o <= x"3C0012AC";
      when 6904 => data_o <= x"00002148";
      when 6905 => data_o <= x"00006BCC";
      when 6906 => data_o <= x"69645FC6";
      when 6907 => data_o <= x"FF524973";
      when 6908 => data_o <= x"0FFF000F";
      when 6909 => data_o <= x"4C0012AC";
      when 6910 => data_o <= x"000021BC";
      when 6911 => data_o <= x"00006BE4";
      when 6912 => data_o <= x"736964C5";
      when 6913 => data_o <= x"FFFF5249";
      when 6914 => data_o <= x"0FFF0013";
      when 6915 => data_o <= x"580012AC";
      when 6916 => data_o <= x"000021F8";
      when 6917 => data_o <= x"00006BFC";
      when 6918 => data_o <= x"61645FC5";
      when 6919 => data_o <= x"FFFF6D73";
      when 6920 => data_o <= x"0FFF0009";
      when 6921 => data_o <= x"610012AC";
      when 6922 => data_o <= x"00002244";
      when 6923 => data_o <= x"00006C14";
      when 6924 => data_o <= x"666564C6";
      when 6925 => data_o <= x"FF3F7265";
      when 6926 => data_o <= x"0FFF0015";
      when 6927 => data_o <= x"680012AC";
      when 6928 => data_o <= x"00002268";
      when 6929 => data_o <= x"00006C2C";
      when 6930 => data_o <= x"736164C4";
      when 6931 => data_o <= x"FFFFFF6D";
      when 6932 => data_o <= x"0FFF002D";
      when 6933 => data_o <= x"740012AC";
      when 6934 => data_o <= x"000022BC";
      when 6935 => data_o <= x"00006C44";
      when 6936 => data_o <= x"656573C3";
      when 6937 => data_o <= x"0FFF0018";
      when 6938 => data_o <= x"860012AC";
      when 6939 => data_o <= x"00002370";
      when 6940 => data_o <= x"00006C5C";
      when 6941 => data_o <= x"636F6CC3";
      when 6942 => data_o <= x"00006CF8";
      when 6943 => data_o <= x"2F2E2E15";
      when 6944 => data_o <= x"662F2E2E";
      when 6945 => data_o <= x"6874726F";
      when 6946 => data_o <= x"726F632F";
      when 6947 => data_o <= x"74786565";
      when 6948 => data_o <= x"FFFF662E";
      when 6949 => data_o <= x"10FF0014";
      when 6950 => data_o <= x"0E0012AC";
      when 6951 => data_o <= x"000023D0";
      when 6952 => data_o <= x"00006C70";
      when 6953 => data_o <= x"756E75C6";
      when 6954 => data_o <= x"FF646573";
      when 6955 => data_o <= x"10FF0005";
      when 6956 => data_o <= x"170012AC";
      when 6957 => data_o <= x"00002420";
      when 6958 => data_o <= x"00006CA0";
      when 6959 => data_o <= x"6C6F72C4";
      when 6960 => data_o <= x"FFFFFF6C";
      when 6961 => data_o <= x"10FF0002";
      when 6962 => data_o <= x"1F0012A4";
      when 6963 => data_o <= x"00002434";
      when 6964 => data_o <= x"00006CB8";
      when 6965 => data_o <= x"6F635BC9";
      when 6966 => data_o <= x"6C69706D";
      when 6967 => data_o <= x"FFFF5D65";
      when 6968 => data_o <= x"10FF0006";
      when 6969 => data_o <= x"220012AC";
      when 6970 => data_o <= x"0000243C";
      when 6971 => data_o <= x"00006CD0";
      when 6972 => data_o <= x"4C4F48C5";
      when 6973 => data_o <= x"FFFF5344";
      when 6974 => data_o <= x"00006D4C";
      when 6975 => data_o <= x"2F2E2E16";
      when 6976 => data_o <= x"662F2E2E";
      when 6977 => data_o <= x"6874726F";
      when 6978 => data_o <= x"6F6F742F";
      when 6979 => data_o <= x"7865736C";
      when 6980 => data_o <= x"FF662E74";
      when 6981 => data_o <= x"11FF0003";
      when 6982 => data_o <= x"030012A4";
      when 6983 => data_o <= x"00002454";
      when 6984 => data_o <= x"00006CEC";
      when 6985 => data_o <= x"65645BC9";
      when 6986 => data_o <= x"656E6966";
      when 6987 => data_o <= x"FFFF5D64";
      when 6988 => data_o <= x"11FF0002";
      when 6989 => data_o <= x"050012A4";
      when 6990 => data_o <= x"00002460";
      when 6991 => data_o <= x"00006D20";
      when 6992 => data_o <= x"6E755BCB";
      when 6993 => data_o <= x"69666564";
      when 6994 => data_o <= x"5D64656E";
      when 6995 => data_o <= x"00006DCC";
      when 6996 => data_o <= x"2F2E2E14";
      when 6997 => data_o <= x"662F2E2E";
      when 6998 => data_o <= x"6874726F";
      when 6999 => data_o <= x"7274732F";
      when 7000 => data_o <= x"2E676E69";
      when 7001 => data_o <= x"FFFFFF66";
      when 7002 => data_o <= x"12FF0012";
      when 7003 => data_o <= x"050012AC";
      when 7004 => data_o <= x"00002468";
      when 7005 => data_o <= x"00006D3C";
      when 7006 => data_o <= x"6D6F63C7";
      when 7007 => data_o <= x"65726170";
      when 7008 => data_o <= x"12FF0002";
      when 7009 => data_o <= x"150012AC";
      when 7010 => data_o <= x"000024B0";
      when 7011 => data_o <= x"00006D74";
      when 7012 => data_o <= x"616C62C5";
      when 7013 => data_o <= x"FFFF6B6E";
      when 7014 => data_o <= x"12FF0007";
      when 7015 => data_o <= x"170012AC";
      when 7016 => data_o <= x"000024B8";
      when 7017 => data_o <= x"00006D8C";
      when 7018 => data_o <= x"72742DC9";
      when 7019 => data_o <= x"696C6961";
      when 7020 => data_o <= x"FFFF676E";
      when 7021 => data_o <= x"12FF0017";
      when 7022 => data_o <= x"210012AC";
      when 7023 => data_o <= x"000024D4";
      when 7024 => data_o <= x"00006DA4";
      when 7025 => data_o <= x"616573C6";
      when 7026 => data_o <= x"FF686372";
      when 7027 => data_o <= x"00007098";
      when 7028 => data_o <= x"2F2E2E14";
      when 7029 => data_o <= x"662F2E2E";
      when 7030 => data_o <= x"6874726F";
      when 7031 => data_o <= x"756F642F";
      when 7032 => data_o <= x"2E656C62";
      when 7033 => data_o <= x"FFFFFF66";
      when 7034 => data_o <= x"13FF0001";
      when 7035 => data_o <= x"030012A8";
      when 7036 => data_o <= x"00002530";
      when 7037 => data_o <= x"00006DC0";
      when 7038 => data_o <= x"733E64C3";
      when 7039 => data_o <= x"13FF0004";
      when 7040 => data_o <= x"040012AC";
      when 7041 => data_o <= x"00002534";
      when 7042 => data_o <= x"00006DF4";
      when 7043 => data_o <= x"6F7232C4";
      when 7044 => data_o <= x"FFFFFF74";
      when 7045 => data_o <= x"13FF0002";
      when 7046 => data_o <= x"050012AC";
      when 7047 => data_o <= x"00002544";
      when 7048 => data_o <= x"00006E08";
      when 7049 => data_o <= x"72322DC5";
      when 7050 => data_o <= x"FFFF746F";
      when 7051 => data_o <= x"13FF0002";
      when 7052 => data_o <= x"060012AC";
      when 7053 => data_o <= x"0000254C";
      when 7054 => data_o <= x"00006E20";
      when 7055 => data_o <= x"696E32C4";
      when 7056 => data_o <= x"FFFFFF70";
      when 7057 => data_o <= x"13FF0002";
      when 7058 => data_o <= x"070012AC";
      when 7059 => data_o <= x"00002554";
      when 7060 => data_o <= x"00006E38";
      when 7061 => data_o <= x"757432C5";
      when 7062 => data_o <= x"FFFF6B63";
      when 7063 => data_o <= x"13FF0002";
      when 7064 => data_o <= x"080012AC";
      when 7065 => data_o <= x"0000255C";
      when 7066 => data_o <= x"00006E50";
      when 7067 => data_o <= x"FF2D64C2";
      when 7068 => data_o <= x"13FF0002";
      when 7069 => data_o <= x"090012AC";
      when 7070 => data_o <= x"00002564";
      when 7071 => data_o <= x"00006E68";
      when 7072 => data_o <= x"FF3C64C2";
      when 7073 => data_o <= x"13FF0002";
      when 7074 => data_o <= x"0A0012AC";
      when 7075 => data_o <= x"0000256C";
      when 7076 => data_o <= x"00006E7C";
      when 7077 => data_o <= x"FF3D64C2";
      when 7078 => data_o <= x"13FF0002";
      when 7079 => data_o <= x"0B0012A8";
      when 7080 => data_o <= x"00002574";
      when 7081 => data_o <= x"00006E90";
      when 7082 => data_o <= x"3D3064C3";
      when 7083 => data_o <= x"13FF0001";
      when 7084 => data_o <= x"0C0012A8";
      when 7085 => data_o <= x"0000257C";
      when 7086 => data_o <= x"00006EA4";
      when 7087 => data_o <= x"3C3064C3";
      when 7088 => data_o <= x"13FF0001";
      when 7089 => data_o <= x"0D0012AC";
      when 7090 => data_o <= x"00002580";
      when 7091 => data_o <= x"00006EB8";
      when 7092 => data_o <= x"2A3264C3";
      when 7093 => data_o <= x"13FF0007";
      when 7094 => data_o <= x"0F0012AC";
      when 7095 => data_o <= x"00002584";
      when 7096 => data_o <= x"00006ECC";
      when 7097 => data_o <= x"2F3264C3";
      when 7098 => data_o <= x"13FF0002";
      when 7099 => data_o <= x"150012A4";
      when 7100 => data_o <= x"000025A0";
      when 7101 => data_o <= x"00006EE0";
      when 7102 => data_o <= x"696C32C8";
      when 7103 => data_o <= x"61726574";
      when 7104 => data_o <= x"FFFFFF6C";
      when 7105 => data_o <= x"13FF0003";
      when 7106 => data_o <= x"1A0012AC";
      when 7107 => data_o <= x"000025A8";
      when 7108 => data_o <= x"00006EF4";
      when 7109 => data_o <= x"617632C9";
      when 7110 => data_o <= x"62616972";
      when 7111 => data_o <= x"FFFF656C";
      when 7112 => data_o <= x"13FF0005";
      when 7113 => data_o <= x"1E0012AC";
      when 7114 => data_o <= x"000025B4";
      when 7115 => data_o <= x"00006F10";
      when 7116 => data_o <= x"6F6332C9";
      when 7117 => data_o <= x"6174736E";
      when 7118 => data_o <= x"FFFF746E";
      when 7119 => data_o <= x"13FF0006";
      when 7120 => data_o <= x"220012AC";
      when 7121 => data_o <= x"000025C8";
      when 7122 => data_o <= x"00006F2C";
      when 7123 => data_o <= x"FF3C64C2";
      when 7124 => data_o <= x"13FF0006";
      when 7125 => data_o <= x"250012AC";
      when 7126 => data_o <= x"000025E0";
      when 7127 => data_o <= x"00006F48";
      when 7128 => data_o <= x"3C7564C3";
      when 7129 => data_o <= x"13FF0006";
      when 7130 => data_o <= x"280012AC";
      when 7131 => data_o <= x"000025F8";
      when 7132 => data_o <= x"00006F5C";
      when 7133 => data_o <= x"616D64C4";
      when 7134 => data_o <= x"FFFFFF78";
      when 7135 => data_o <= x"13FF0007";
      when 7136 => data_o <= x"2B0012AC";
      when 7137 => data_o <= x"00002610";
      when 7138 => data_o <= x"00006F70";
      when 7139 => data_o <= x"696D64C4";
      when 7140 => data_o <= x"FFFFFF6E";
      when 7141 => data_o <= x"13FF0002";
      when 7142 => data_o <= x"2F0012AC";
      when 7143 => data_o <= x"0000262C";
      when 7144 => data_o <= x"00006F88";
      when 7145 => data_o <= x"FF2B6DC2";
      when 7146 => data_o <= x"13FF0008";
      when 7147 => data_o <= x"310012AC";
      when 7148 => data_o <= x"00002634";
      when 7149 => data_o <= x"00006FA0";
      when 7150 => data_o <= x"FF2A6DC2";
      when 7151 => data_o <= x"13FF0006";
      when 7152 => data_o <= x"3A0012AC";
      when 7153 => data_o <= x"00002654";
      when 7154 => data_o <= x"00006FB4";
      when 7155 => data_o <= x"656E74C7";
      when 7156 => data_o <= x"65746167";
      when 7157 => data_o <= x"13FF000D";
      when 7158 => data_o <= x"3E0012AC";
      when 7159 => data_o <= x"0000266C";
      when 7160 => data_o <= x"00006FC8";
      when 7161 => data_o <= x"FF2A74C2";
      when 7162 => data_o <= x"13FF000B";
      when 7163 => data_o <= x"480012AC";
      when 7164 => data_o <= x"000026A0";
      when 7165 => data_o <= x"00006FE0";
      when 7166 => data_o <= x"FF2F74C2";
      when 7167 => data_o <= x"13FF0002";
      when 7168 => data_o <= x"520012AC";
      when 7169 => data_o <= x"000026CC";
      when 7170 => data_o <= x"00006FF4";
      when 7171 => data_o <= x"2F2A6DC3";
      when 7172 => data_o <= x"00FF000B";
      when 7173 => data_o <= x"430012AC";
      when 7174 => data_o <= x"000026D4";
      when 7175 => data_o <= x"00007008";
      when 7176 => data_o <= x"69616DC4";
      when 7177 => data_o <= x"FFFFFF6E";
      when 7178 => data_o <= x"00FF000B";
      when 7179 => data_o <= x"480012AC";
      when 7180 => data_o <= x"00002700";
      when 7181 => data_o <= x"0000701C";
      when 7182 => data_o <= x"424946C3";
      when 7183 => data_o <= x"00FF0004";
      when 7184 => data_o <= x"4E0012AC";
      when 7185 => data_o <= x"0000272C";
      when 7186 => data_o <= x"00007034";
      when 7187 => data_o <= x"6D6F74C4";
      when 7188 => data_o <= x"FFFFFF73";
      when 7189 => data_o <= x"00FF0019";
      when 7190 => data_o <= x"520012AC";
      when 7191 => data_o <= x"0000273C";
      when 7192 => data_o <= x"00007048";
      when 7193 => data_o <= x"6E6562C5";
      when 7194 => data_o <= x"FFFF6863";
      when 7195 => data_o <= x"00FF0004";
      when 7196 => data_o <= x"590012AC";
      when 7197 => data_o <= x"000027A0";
      when 7198 => data_o <= x"00007060";
      when 7199 => data_o <= x"316666C4";
      when 7200 => data_o <= x"FFFFFF64";
      when 7201 => data_o <= x"00FF0002";
      when 7202 => data_o <= x"5E0012AC";
      when 7203 => data_o <= x"000027B0";
      when 7204 => data_o <= x"00007078";
      when 7205 => data_o <= x"316666C3";
      when 7206 => data_o <= x"FFFFFFFF";
      when 7207 => data_o <= x"2F2E2E11";
      when 7208 => data_o <= x"662F2E2E";
      when 7209 => data_o <= x"6874726F";
      when 7210 => data_o <= x"646E652F";
      when 7211 => data_o <= x"FFFF662E";
      when 7212 => data_o <= x"000027B8";
      when 7213 => data_o <= x"14FFFFFF";
      when 7214 => data_o <= x"040012BC";
      when 7215 => data_o <= x"000012B8";
      when 7216 => data_o <= x"00007090";
      when 7217 => data_o <= x"6164490A";
      when 7218 => data_o <= x"61546174";
      when 7219 => data_o <= x"FF656C62";
      when 7220 => data_o <= x"14FF0017";
      when 7221 => data_o <= x"070012AC";
      when 7222 => data_o <= x"00002844";
      when 7223 => data_o <= x"000070C0";
      when 7224 => data_o <= x"696E694A";
      when 7225 => data_o <= x"6C616974";
      when 7226 => data_o <= x"FF657A69";
      when others => data_o <= x"00000000";
    end case;
  end if;
end process;

END ARCHITECTURE RTL;
