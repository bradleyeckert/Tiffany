library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

-- Single-port synchronous-read ROM

ENTITY ROM32 IS
generic (
  Size:  integer := 10                          -- log2 (cells)
);
port (
  clk:    in  std_logic;                        -- System clock
  addr:   in  std_logic_vector(Size-1 downto 0);
  data_o: out std_logic_vector(31 downto 0)     -- read data
);
END ROM32;

ARCHITECTURE RTL OF ROM32 IS
signal address: integer range 0 to 2**Size-1;
begin
address <= to_integer(unsigned(addr));

process (address) begin
  if rising_edge(clk) then
    case address is
      when   0 => data_o <= x"5400028A";
      when   1 => data_o <= x"5400028D";
      when   2 => data_o <= x"57FFFFFF";
      when   3 => data_o <= x"D090C220";
      when   4 => data_o <= x"9FB08800";
      when   5 => data_o <= x"3FB08800";
      when   6 => data_o <= x"5FB08800";
      when   7 => data_o <= x"05FB8318";
      when   8 => data_o <= x"9FB08800";
      when   9 => data_o <= x"05FD8318";
      when  10 => data_o <= x"3FB08800";
      when  11 => data_o <= x"D0908800";
      when  12 => data_o <= x"D09D0220";
      when  13 => data_o <= x"D21D0220";
      when  14 => data_o <= x"10408800";
      when  15 => data_o <= x"7FC1BC08";
      when  16 => data_o <= x"F1FF0608";
      when  17 => data_o <= x"F3908800";
      when  18 => data_o <= x"F3B08800";
      when  19 => data_o <= x"F06F1FF0";
      when  20 => data_o <= x"7DF08800";
      when  21 => data_o <= x"186F06F0";
      when  22 => data_o <= x"7FC08800";
      when  23 => data_o <= x"186FBC7C";
      when  24 => data_o <= x"F3EF1F08";
      when  25 => data_o <= x"EFB08800";
      when  26 => data_o <= x"E7908800";
      when  27 => data_o <= x"7FC1BC7C";
      when  28 => data_o <= x"7FC1BC1A";
      when  29 => data_o <= x"7DFE7918";
      when  30 => data_o <= x"1950001B";
      when  31 => data_o <= x"EFBEC220";
      when  32 => data_o <= x"07A08800";
      when  33 => data_o <= x"04220000";
      when  34 => data_o <= x"07005BD2";
      when  35 => data_o <= x"05B08800";
      when  36 => data_o <= x"90220000";
      when  37 => data_o <= x"6E408800";
      when  38 => data_o <= x"6E490220";
      when  39 => data_o <= x"92408800";
      when  40 => data_o <= x"D09B0220";
      when  41 => data_o <= x"24927D03";
      when  42 => data_o <= x"D1308800";
      when  43 => data_o <= x"9BCBBC08";
      when  44 => data_o <= x"9E7EC220";
      when  45 => data_o <= x"C3424800";
      when  46 => data_o <= x"08800000";
      when  47 => data_o <= x"D3CD13D2";
      when  48 => data_o <= x"7C220000";
      when  49 => data_o <= x"7DFF060C";
      when  50 => data_o <= x"F068C220";
      when  51 => data_o <= x"D1FD0918";
      when  52 => data_o <= x"E64C3B26";
      when  53 => data_o <= x"EC220000";
      when  54 => data_o <= x"C1500033";
      when  55 => data_o <= x"08800000";
      when  56 => data_o <= x"38220000";
      when  57 => data_o <= x"F4000004";
      when  58 => data_o <= x"66E08800";
      when  59 => data_o <= x"F4000008";
      when  60 => data_o <= x"66E08800";
      when  61 => data_o <= x"F400000C";
      when  62 => data_o <= x"A6EF4008";
      when  63 => data_o <= x"67424350";
      when  64 => data_o <= x"50220000";
      when  65 => data_o <= x"044119B8";
      when  66 => data_o <= x"F3B08800";
      when  67 => data_o <= x"F400000A";
      when  68 => data_o <= x"F4000DE7";
      when  69 => data_o <= x"D27EC220";
      when  70 => data_o <= x"F4000010";
      when  71 => data_o <= x"F4000DE7";
      when  72 => data_o <= x"D27EC220";
      when  73 => data_o <= x"B8800000";
      when  74 => data_o <= x"F4FFFFFF";
      when  75 => data_o <= x"4C220000";
      when  76 => data_o <= x"E79D0320";
      when  77 => data_o <= x"C3BEFB08";
      when  78 => data_o <= x"EFCD0918";
      when  79 => data_o <= x"87C7FC7C";
      when  80 => data_o <= x"7C220000";
      when  81 => data_o <= x"186246E4";
      when  82 => data_o <= x"E4320000";
      when  83 => data_o <= x"C3B7DF7E";
      when  84 => data_o <= x"EFBEE17E";
      when  85 => data_o <= x"1BC1B90C";
      when  86 => data_o <= x"FB90FC7C";
      when  87 => data_o <= x"F2C6C800";
      when  88 => data_o <= x"C3B7C220";
      when  89 => data_o <= x"EC6EC6EC";
      when  90 => data_o <= x"85F08800";
      when  91 => data_o <= x"F400000C";
      when  92 => data_o <= x"46E08800";
      when  93 => data_o <= x"186EC6EC";
      when  94 => data_o <= x"7C220000";
      when  95 => data_o <= x"E796E420";
      when  96 => data_o <= x"EBB08800";
      when  97 => data_o <= x"EFB1A17E";
      when  98 => data_o <= x"186D09D0";
      when  99 => data_o <= x"C3B7C220";
      when 100 => data_o <= x"7E17C220";
      when 101 => data_o <= x"181383F7";
      when 102 => data_o <= x"05F0C6D0";
      when 103 => data_o <= x"4DF08800";
      when 104 => data_o <= x"E796EC20";
      when 105 => data_o <= x"EB4243B2";
      when 106 => data_o <= x"F3BB0220";
      when 107 => data_o <= x"F1500068";
      when 108 => data_o <= x"E796EC20";
      when 109 => data_o <= x"EB4243B2";
      when 110 => data_o <= x"EEC08800";
      when 111 => data_o <= x"F150006C";
      when 112 => data_o <= x"D09D0800";
      when 113 => data_o <= x"C1500075";
      when 114 => data_o <= x"D09F1FF0";
      when 115 => data_o <= x"9869DFA0";
      when 116 => data_o <= x"1BBEFB08";
      when 117 => data_o <= x"EFBEC220";
      when 118 => data_o <= x"D09D0800";
      when 119 => data_o <= x"C150007B";
      when 120 => data_o <= x"D09F1FF0";
      when 121 => data_o <= x"3863DFA0";
      when 122 => data_o <= x"1BBEFB08";
      when 123 => data_o <= x"EFBEC220";
      when 124 => data_o <= x"D09D0800";
      when 125 => data_o <= x"C1500085";
      when 126 => data_o <= x"2417C3F0";
      when 127 => data_o <= x"F83F06D0";
      when 128 => data_o <= x"24800000";
      when 129 => data_o <= x"7F4274F0";
      when 130 => data_o <= x"D09D3CE4";
      when 131 => data_o <= x"DB93FB18";
      when 132 => data_o <= x"27054081";
      when 133 => data_o <= x"EFBEC220";
      when 134 => data_o <= x"7F9E5D68";
      when 135 => data_o <= x"E950008A";
      when 136 => data_o <= x"19D0007C";
      when 137 => data_o <= x"5400008B";
      when 138 => data_o <= x"19D00076";
      when 139 => data_o <= x"08800000";
      when 140 => data_o <= x"E7A54091";
      when 141 => data_o <= x"F34249F0";
      when 142 => data_o <= x"7FC20000";
      when 143 => data_o <= x"FBC3E818";
      when 144 => data_o <= x"EFBEC220";
      when 145 => data_o <= x"EFBEC220";
      when 146 => data_o <= x"F4000000";
      when 147 => data_o <= x"5400008C";
      when 148 => data_o <= x"D09D30EE";
      when 149 => data_o <= x"F400003F";
      when 150 => data_o <= x"4F427C20";
      when 151 => data_o <= x"128F3B08";
      when 152 => data_o <= x"08800000";
      when 153 => data_o <= x"D09D30EE";
      when 154 => data_o <= x"F400003F";
      when 155 => data_o <= x"4F427C20";
      when 156 => data_o <= x"728F3B08";
      when 157 => data_o <= x"08800000";
      when 158 => data_o <= x"0416FD1F";
      when 159 => data_o <= x"D0800000";
      when 160 => data_o <= x"7C47CC20";
      when 161 => data_o <= x"E391837C";
      when 162 => data_o <= x"E0920000";
      when 163 => data_o <= x"18624800";
      when 164 => data_o <= x"C15000A0";
      when 165 => data_o <= x"EDF7FB18";
      when 166 => data_o <= x"1BC08800";
      when 167 => data_o <= x"E79D090C";
      when 168 => data_o <= x"EF8540B7";
      when 169 => data_o <= x"F400001F";
      when 170 => data_o <= x"D1C10800";
      when 171 => data_o <= x"7DF7CC18";
      when 172 => data_o <= x"338540B2";
      when 173 => data_o <= x"07ED090C";
      when 174 => data_o <= x"EC800000";
      when 175 => data_o <= x"E3ED090C";
      when 176 => data_o <= x"04CD14EC";
      when 177 => data_o <= x"540000B4";
      when 178 => data_o <= x"FB4243F4";
      when 179 => data_o <= x"13B20000";
      when 180 => data_o <= x"18624800";
      when 181 => data_o <= x"C15000AB";
      when 182 => data_o <= x"EFBF0CD2";
      when 183 => data_o <= x"EFBEFD00";
      when 184 => data_o <= x"D0108800";
      when 185 => data_o <= x"E796DFE4";
      when 186 => data_o <= x"7DD0002D";
      when 187 => data_o <= x"7DD00036";
      when 188 => data_o <= x"19D000A7";
      when 189 => data_o <= x"F06B0800";
      when 190 => data_o <= x"E95000C0";
      when 191 => data_o <= x"D0920000";
      when 192 => data_o <= x"F06B0800";
      when 193 => data_o <= x"E95000C3";
      when 194 => data_o <= x"D0920000";
      when 195 => data_o <= x"08800000";
      when 196 => data_o <= x"05FE796C";
      when 197 => data_o <= x"7C17DD2D";
      when 198 => data_o <= x"7DD00036";
      when 199 => data_o <= x"19D000A7";
      when 200 => data_o <= x"F06B0800";
      when 201 => data_o <= x"E95000CB";
      when 202 => data_o <= x"D0920000";
      when 203 => data_o <= x"F06B0800";
      when 204 => data_o <= x"E95000D2";
      when 205 => data_o <= x"D09E4800";
      when 206 => data_o <= x"E95000D2";
      when 207 => data_o <= x"F9FF06F0";
      when 208 => data_o <= x"D090FCD0";
      when 209 => data_o <= x"27420000";
      when 210 => data_o <= x"1BB08800";
      when 211 => data_o <= x"06C05F20";
      when 212 => data_o <= x"E95000D7";
      when 213 => data_o <= x"D097DD33";
      when 214 => data_o <= x"18800000";
      when 215 => data_o <= x"7C1B0800";
      when 216 => data_o <= x"E95000DA";
      when 217 => data_o <= x"F8320000";
      when 218 => data_o <= x"19D000A7";
      when 219 => data_o <= x"1BA540DD";
      when 220 => data_o <= x"F3427C20";
      when 221 => data_o <= x"08800000";
      when 222 => data_o <= x"E6CF15D3";
      when 223 => data_o <= x"740000DE";
      when 224 => data_o <= x"EC220000";
      when 225 => data_o <= x"740000DE";
      when 226 => data_o <= x"F3B08800";
      when 227 => data_o <= x"E797406C";
      when 228 => data_o <= x"EBC20000";
      when 229 => data_o <= x"EC220000";
      when 230 => data_o <= x"E79F1D6C";
      when 231 => data_o <= x"EBC20000";
      when 232 => data_o <= x"EC220000";
      when 233 => data_o <= x"E7974068";
      when 234 => data_o <= x"EBC20000";
      when 235 => data_o <= x"EC220000";
      when 236 => data_o <= x"E79F1D68";
      when 237 => data_o <= x"EBC20000";
      when 238 => data_o <= x"EC220000";
      when 239 => data_o <= x"7FCF83F0";
      when 240 => data_o <= x"1B424308";
      when 241 => data_o <= x"E742437C";
      when 242 => data_o <= x"D090C620";
      when 243 => data_o <= x"54000068";
      when 244 => data_o <= x"7400009E";
      when 245 => data_o <= x"EC220000";
      when 246 => data_o <= x"E796EC7C";
      when 247 => data_o <= x"7400002D";
      when 248 => data_o <= x"F1D0002D";
      when 249 => data_o <= x"7400009E";
      when 250 => data_o <= x"1BA540FC";
      when 251 => data_o <= x"74000033";
      when 252 => data_o <= x"08800000";
      when 253 => data_o <= x"7DD000F6";
      when 254 => data_o <= x"195000D3";
      when 255 => data_o <= x"740000FD";
      when 256 => data_o <= x"F3B08800";
      when 257 => data_o <= x"34000006";
      when 258 => data_o <= x"08800000";
      when 259 => data_o <= x"F3D00000";
      when 260 => data_o <= x"D1F20000";
      when 261 => data_o <= x"E7A5410F";
      when 262 => data_o <= x"F34274F0";
      when 263 => data_o <= x"3866FD07";
      when 264 => data_o <= x"D0800000";
      when 265 => data_o <= x"25F07D01";
      when 266 => data_o <= x"4F427DED";
      when 267 => data_o <= x"94B88320";
      when 268 => data_o <= x"4FC71B18";
      when 269 => data_o <= x"C1500109";
      when 270 => data_o <= x"EDF54105";
      when 271 => data_o <= x"EFB1B408";
      when 272 => data_o <= x"E5FF4004";
      when 273 => data_o <= x"65FF4DEB";
      when 274 => data_o <= x"D2E7FD00";
      when 275 => data_o <= x"47D00DEB";
      when 276 => data_o <= x"D27EDD30";
      when 277 => data_o <= x"1BD00DEB";
      when 278 => data_o <= x"D27EC6EC";
      when 279 => data_o <= x"1816C220";
      when 280 => data_o <= x"07AEC220";
      when 281 => data_o <= x"F4000DEB";
      when 282 => data_o <= x"D2EBC620";
      when 283 => data_o <= x"F4000DEB";
      when 284 => data_o <= x"D27EC6F0";
      when 285 => data_o <= x"7F7EFCEC";
      when 286 => data_o <= x"186F0220";
      when 287 => data_o <= x"08800000";
      when 288 => data_o <= x"04D00004";
      when 289 => data_o <= x"08800000";
      when 290 => data_o <= x"F400000A";
      when 291 => data_o <= x"740000F4";
      when 292 => data_o <= x"74000120";
      when 293 => data_o <= x"0C800000";
      when 294 => data_o <= x"7400011F";
      when 295 => data_o <= x"05D00120";
      when 296 => data_o <= x"7400006C";
      when 297 => data_o <= x"E9500126";
      when 298 => data_o <= x"EC220000";
      when 299 => data_o <= x"7400011F";
      when 300 => data_o <= x"04D00003";
      when 301 => data_o <= x"E950012B";
      when 302 => data_o <= x"34000002";
      when 303 => data_o <= x"EC220000";
      when 304 => data_o <= x"5400016F";
      when 305 => data_o <= x"39500130";
      when 306 => data_o <= x"040A0D02";
      when 307 => data_o <= x"4A325B1B";
      when 308 => data_o <= x"F40004C8";
      when 309 => data_o <= x"54000131";
      when 310 => data_o <= x"F40004CB";
      when 311 => data_o <= x"54000131";
      when 312 => data_o <= x"04D00000";
      when 313 => data_o <= x"5400011F";
      when 314 => data_o <= x"74000138";
      when 315 => data_o <= x"E950013A";
      when 316 => data_o <= x"04D00001";
      when 317 => data_o <= x"08800000";
      when 318 => data_o <= x"000004AC";
      when 319 => data_o <= x"000004D0";
      when 320 => data_o <= x"000004D8";
      when 321 => data_o <= x"000004E0";
      when 322 => data_o <= x"000004E8";
      when 323 => data_o <= x"F40004F8";
      when 324 => data_o <= x"F4000DCF";
      when 325 => data_o <= x"D27EC220";
      when 326 => data_o <= x"104F4DCF";
      when 327 => data_o <= x"D2E0EE7E";
      when 328 => data_o <= x"F4000000";
      when 329 => data_o <= x"54000146";
      when 330 => data_o <= x"F4000001";
      when 331 => data_o <= x"54000146";
      when 332 => data_o <= x"F4000002";
      when 333 => data_o <= x"54000146";
      when 334 => data_o <= x"F4000003";
      when 335 => data_o <= x"54000146";
      when 336 => data_o <= x"F4000004";
      when 337 => data_o <= x"54000146";
      when 338 => data_o <= x"E5FD09D0";
      when 339 => data_o <= x"F09F06DA";
      when 340 => data_o <= x"F4000006";
      when 341 => data_o <= x"74000094";
      when 342 => data_o <= x"7DD00152";
      when 343 => data_o <= x"F400003F";
      when 344 => data_o <= x"4C60C220";
      when 345 => data_o <= x"74000152";
      when 346 => data_o <= x"07D000C0";
      when 347 => data_o <= x"4FD00080";
      when 348 => data_o <= x"6E420000";
      when 349 => data_o <= x"E950015F";
      when 350 => data_o <= x"ED500159";
      when 351 => data_o <= x"07D00080";
      when 352 => data_o <= x"4FA5416E";
      when 353 => data_o <= x"07D00020";
      when 354 => data_o <= x"4FA5416C";
      when 355 => data_o <= x"07D00010";
      when 356 => data_o <= x"4FA54169";
      when 357 => data_o <= x"F4000007";
      when 358 => data_o <= x"4DD00154";
      when 359 => data_o <= x"74000154";
      when 360 => data_o <= x"54000154";
      when 361 => data_o <= x"F400000F";
      when 362 => data_o <= x"4DD00154";
      when 363 => data_o <= x"54000154";
      when 364 => data_o <= x"F400001F";
      when 365 => data_o <= x"4D500154";
      when 366 => data_o <= x"08800000";
      when 367 => data_o <= x"074274B0";
      when 368 => data_o <= x"D3A54174";
      when 369 => data_o <= x"74000159";
      when 370 => data_o <= x"74000148";
      when 371 => data_o <= x"5400016F";
      when 372 => data_o <= x"EFB08800";
      when 373 => data_o <= x"F4000020";
      when 374 => data_o <= x"54000148";
      when 375 => data_o <= x"C3B08800";
      when 376 => data_o <= x"74000175";
      when 377 => data_o <= x"D09D0800";
      when 378 => data_o <= x"54000177";
      when 379 => data_o <= x"08800000";
      when 380 => data_o <= x"F4000009";
      when 381 => data_o <= x"E5D0006C";
      when 382 => data_o <= x"F4000007";
      when 383 => data_o <= x"4C3F4030";
      when 384 => data_o <= x"0C220000";
      when 385 => data_o <= x"F4000CCB";
      when 386 => data_o <= x"D3D00D97";
      when 387 => data_o <= x"D27EC220";
      when 388 => data_o <= x"F4000D97";
      when 389 => data_o <= x"D2ED09D1";
      when 390 => data_o <= x"F4000D97";
      when 391 => data_o <= x"D27ECFEE";
      when 392 => data_o <= x"F4000000";
      when 393 => data_o <= x"F4000DE7";
      when 394 => data_o <= x"D2E740A7";
      when 395 => data_o <= x"7FD00DE7";
      when 396 => data_o <= x"D2E740A7";
      when 397 => data_o <= x"F1D0017C";
      when 398 => data_o <= x"74000184";
      when 399 => data_o <= x"18220000";
      when 400 => data_o <= x"74000188";
      when 401 => data_o <= x"E797402F";
      when 402 => data_o <= x"93A54190";
      when 403 => data_o <= x"08800000";
      when 404 => data_o <= x"B3A54197";
      when 405 => data_o <= x"F400002D";
      when 406 => data_o <= x"74000184";
      when 407 => data_o <= x"08800000";
      when 408 => data_o <= x"EFBF4D97";
      when 409 => data_o <= x"D2EF4CCB";
      when 410 => data_o <= x"D39D090E";
      when 411 => data_o <= x"E7424320";
      when 412 => data_o <= x"74000177";
      when 413 => data_o <= x"54000130";
      when 414 => data_o <= x"7C17DD36";
      when 415 => data_o <= x"74000181";
      when 416 => data_o <= x"74000190";
      when 417 => data_o <= x"19D00194";
      when 418 => data_o <= x"74000198";
      when 419 => data_o <= x"1950019B";
      when 420 => data_o <= x"F4000000";
      when 421 => data_o <= x"F150019E";
      when 422 => data_o <= x"7DD00022";
      when 423 => data_o <= x"1950019E";
      when 424 => data_o <= x"F4000000";
      when 425 => data_o <= x"7400019E";
      when 426 => data_o <= x"54000175";
      when 427 => data_o <= x"F4000000";
      when 428 => data_o <= x"540001A8";
      when 429 => data_o <= x"F4000DE7";
      when 430 => data_o <= x"D2EF400A";
      when 431 => data_o <= x"6FA541B1";
      when 432 => data_o <= x"540001AB";
      when 433 => data_o <= x"74000022";
      when 434 => data_o <= x"540001A8";
      when 435 => data_o <= x"B95001AD";
      when 436 => data_o <= x"74000181";
      when 437 => data_o <= x"D0920000";
      when 438 => data_o <= x"7DD00188";
      when 439 => data_o <= x"18920000";
      when 440 => data_o <= x"C15001B6";
      when 441 => data_o <= x"EDD00190";
      when 442 => data_o <= x"54000198";
      when 443 => data_o <= x"F4000DE7";
      when 444 => data_o <= x"D2E7DD46";
      when 445 => data_o <= x"F4000000";
      when 446 => data_o <= x"F1D001B4";
      when 447 => data_o <= x"1BD00DE7";
      when 448 => data_o <= x"D27EC800";
      when 449 => data_o <= x"74000130";
      when 450 => data_o <= x"54000175";
      when 451 => data_o <= x"7C10460C";
      when 452 => data_o <= x"7C800000";
      when 453 => data_o <= x"07E6C800";
      when 454 => data_o <= x"E95001E7";
      when 455 => data_o <= x"7400011F";
      when 456 => data_o <= x"7400014E";
      when 457 => data_o <= x"E95001C7";
      when 458 => data_o <= x"74000150";
      when 459 => data_o <= x"07D0000D";
      when 460 => data_o <= x"6E420000";
      when 461 => data_o <= x"E95001D0";
      when 462 => data_o <= x"EC6EFCD0";
      when 463 => data_o <= x"24308800";
      when 464 => data_o <= x"07D00008";
      when 465 => data_o <= x"6E420000";
      when 466 => data_o <= x"E95001DC";
      when 467 => data_o <= x"EF9E5B20";
      when 468 => data_o <= x"E95001DB";
      when 469 => data_o <= x"D09D0800";
      when 470 => data_o <= x"540001D9";
      when 471 => data_o <= x"445B1B07";
      when 472 => data_o <= x"445B1B20";
      when 473 => data_o <= x"F400075C";
      when 474 => data_o <= x"39D00130";
      when 475 => data_o <= x"540001E6";
      when 476 => data_o <= x"07D00020";
      when 477 => data_o <= x"D090C800";
      when 478 => data_o <= x"C15001E5";
      when 479 => data_o <= x"EFD00DB1";
      when 480 => data_o <= x"D3690800";
      when 481 => data_o <= x"E95001E3";
      when 482 => data_o <= x"05D00148";
      when 483 => data_o <= x"F0F20000";
      when 484 => data_o <= x"540001E6";
      when 485 => data_o <= x"EFB20000";
      when 486 => data_o <= x"540001C5";
      when 487 => data_o <= x"1BBF3427";
      when 488 => data_o <= x"08800000";
      when 489 => data_o <= x"9FB08800";
      when 490 => data_o <= x"7F4F40FF";
      when 491 => data_o <= x"4FEF4003";
      when 492 => data_o <= x"4C410420";
      when 493 => data_o <= x"74000094";
      when 494 => data_o <= x"D06F4003";
      when 495 => data_o <= x"D139FB08";
      when 496 => data_o <= x"D0920000";
      when 497 => data_o <= x"7F9DB920";
      when 498 => data_o <= x"740001EA";
      when 499 => data_o <= x"27C27C18";
      when 500 => data_o <= x"270541F1";
      when 501 => data_o <= x"EFBEC220";
      when 502 => data_o <= x"F4000000";
      when 503 => data_o <= x"F4000D9C";
      when 504 => data_o <= x"D0FEC220";
      when 505 => data_o <= x"F4000001";
      when 506 => data_o <= x"F4000D9C";
      when 507 => data_o <= x"D0FEC220";
      when 508 => data_o <= x"F4000D9C";
      when 509 => data_o <= x"D3620000";
      when 510 => data_o <= x"E9500201";
      when 511 => data_o <= x"F4000DDF";
      when 512 => data_o <= x"D0220000";
      when 513 => data_o <= x"F4000DDB";
      when 514 => data_o <= x"D0220000";
      when 515 => data_o <= x"05FB8800";
      when 516 => data_o <= x"740001E9";
      when 517 => data_o <= x"F4000004";
      when 518 => data_o <= x"19500007";
      when 519 => data_o <= x"F4000DDF";
      when 520 => data_o <= x"D1500203";
      when 521 => data_o <= x"F4000DE3";
      when 522 => data_o <= x"D1500203";
      when 523 => data_o <= x"F4000DDB";
      when 524 => data_o <= x"D017EE9C";
      when 525 => data_o <= x"EFD00004";
      when 526 => data_o <= x"19500007";
      when 527 => data_o <= x"F4000D9C";
      when 528 => data_o <= x"D3620000";
      when 529 => data_o <= x"E9500213";
      when 530 => data_o <= x"54000207";
      when 531 => data_o <= x"5400020B";
      when 532 => data_o <= x"05FB8800";
      when 533 => data_o <= x"740001EA";
      when 534 => data_o <= x"FAE2469C";
      when 535 => data_o <= x"EC220000";
      when 536 => data_o <= x"F4000DDF";
      when 537 => data_o <= x"D1500214";
      when 538 => data_o <= x"F4000DE3";
      when 539 => data_o <= x"D1500214";
      when 540 => data_o <= x"F4000DDB";
      when 541 => data_o <= x"D017EE3C";
      when 542 => data_o <= x"EFD00001";
      when 543 => data_o <= x"19500007";
      when 544 => data_o <= x"F4000D9C";
      when 545 => data_o <= x"D3620000";
      when 546 => data_o <= x"E9500224";
      when 547 => data_o <= x"54000218";
      when 548 => data_o <= x"5400021C";
      when 549 => data_o <= x"E7D00DDB";
      when 550 => data_o <= x"D2E6D308";
      when 551 => data_o <= x"F4000DDF";
      when 552 => data_o <= x"D2EF3D00";
      when 553 => data_o <= x"D1D00207";
      when 554 => data_o <= x"06E90800";
      when 555 => data_o <= x"74000225";
      when 556 => data_o <= x"E950022E";
      when 557 => data_o <= x"8550022A";
      when 558 => data_o <= x"04174207";
      when 559 => data_o <= x"06E92420";
      when 560 => data_o <= x"74000225";
      when 561 => data_o <= x"E9500234";
      when 562 => data_o <= x"99D00207";
      when 563 => data_o <= x"5400022F";
      when 564 => data_o <= x"08800000";
      when 565 => data_o <= x"F4000DC7";
      when 566 => data_o <= x"D2EF4DBF";
      when 567 => data_o <= x"D27EC800";
      when 568 => data_o <= x"F4000D97";
      when 569 => data_o <= x"D3D000CC";
      when 570 => data_o <= x"74000092";
      when 571 => data_o <= x"F4000000";
      when 572 => data_o <= x"A4800000";
      when 573 => data_o <= x"74000227";
      when 574 => data_o <= x"7F427E0C";
      when 575 => data_o <= x"514F39F0";
      when 576 => data_o <= x"740001E9";
      when 577 => data_o <= x"1BC90800";
      when 578 => data_o <= x"E950023D";
      when 579 => data_o <= x"EC220000";
      when 580 => data_o <= x"54000249";
      when 581 => data_o <= x"6C65480C";
      when 582 => data_o <= x"57206F6C";
      when 583 => data_o <= x"646C726F";
      when 584 => data_o <= x"FFFFFF21";
      when 585 => data_o <= x"F4000914";
      when 586 => data_o <= x"39D00130";
      when 587 => data_o <= x"7400014A";
      when 588 => data_o <= x"F400000A";
      when 589 => data_o <= x"F4000000";
      when 590 => data_o <= x"F3425F7C";
      when 591 => data_o <= x"F9D001AD";
      when 592 => data_o <= x"74000051";
      when 593 => data_o <= x"5400024F";
      when 594 => data_o <= x"08800000";
      when 595 => data_o <= x"00000003";
      when 596 => data_o <= x"FFFFF204";
      when 597 => data_o <= x"FFFFF200";
      when 598 => data_o <= x"FFFFF1F0";
      when 599 => data_o <= x"FFFFF100";
      when 600 => data_o <= x"00000004";
      when 601 => data_o <= x"FFFFF218";
      when 602 => data_o <= x"0000000A";
      when 603 => data_o <= x"0000A4BC";
      when 604 => data_o <= x"00000970";
      when 605 => data_o <= x"FFFFF338";
      when 606 => data_o <= x"00000006";
      when 607 => data_o <= x"FFFFF22C";
      when 608 => data_o <= x"FFFFF334";
      when 609 => data_o <= x"000004F8";
      when 610 => data_o <= x"00000001";
      when 611 => data_o <= x"0000000C";
      when 612 => data_o <= x"FFFFF26C";
      when 613 => data_o <= x"0000000C";
      when 614 => data_o <= x"00000001";
      when 615 => data_o <= x"FFFFF248";
      when 616 => data_o <= x"001A0001";
      when 617 => data_o <= x"00000001";
      when 618 => data_o <= x"FFFFF250";
      when 619 => data_o <= x"1A000944";
      when 620 => data_o <= x"00000003";
      when 621 => data_o <= x"FFFFF25C";
      when 622 => data_o <= x"0000A480";
      when 623 => data_o <= x"00050003";
      when 624 => data_o <= x"FFFFF334";
      when 625 => data_o <= x"00000001";
      when 626 => data_o <= x"FFFFF334";
      when 627 => data_o <= x"0000A498";
      when 628 => data_o <= x"00000000";
      when 629 => data_o <= x"FFFFF338";
      when 630 => data_o <= x"F400094C";
      when 631 => data_o <= x"9B9E4910";
      when 632 => data_o <= x"103F1FF0";
      when 633 => data_o <= x"18120000";
      when 634 => data_o <= x"E950027D";
      when 635 => data_o <= x"7E619D70";
      when 636 => data_o <= x"54000277";
      when 637 => data_o <= x"1BD00D97";
      when 638 => data_o <= x"D27EC800";
      when 639 => data_o <= x"F4000DFF";
      when 640 => data_o <= x"D3FF4EFF";
      when 641 => data_o <= x"D37F4E13";
      when 642 => data_o <= x"D2FF4D97";
      when 643 => data_o <= x"D2E7C800";
      when 644 => data_o <= x"F4010000";
      when 645 => data_o <= x"F4000DDF";
      when 646 => data_o <= x"D27EC800";
      when 647 => data_o <= x"F4018000";
      when 648 => data_o <= x"F4000DE3";
      when 649 => data_o <= x"D27EC220";
      when 650 => data_o <= x"74000276";
      when 651 => data_o <= x"74000244";
      when 652 => data_o <= x"54000101";
      when 653 => data_o <= x"74000276";
      when 654 => data_o <= x"74000244";
      when 655 => data_o <= x"54000101";
      when others => data_o <= x"00000000";
    end case;
  end if;
end process;

END ARCHITECTURE RTL;
